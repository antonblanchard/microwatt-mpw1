magic
tech sky130A
magscale 1 2
timestamp 1611917162
<< obsli1 >>
rect 1104 2159 582820 701777
<< obsm1 >>
rect 566 2128 582820 701808
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703520
rect 8254 703464 24222 703520
rect 24446 703464 40414 703520
rect 40638 703464 56698 703520
rect 56922 703464 72890 703520
rect 73114 703464 89082 703520
rect 89306 703464 105366 703520
rect 105590 703464 121558 703520
rect 121782 703464 137750 703520
rect 137974 703464 154034 703520
rect 154258 703464 170226 703520
rect 170450 703464 186418 703520
rect 186642 703464 202702 703520
rect 202926 703464 218894 703520
rect 219118 703464 235086 703520
rect 235310 703464 251370 703520
rect 251594 703464 267562 703520
rect 267786 703464 283754 703520
rect 283978 703464 300038 703520
rect 300262 703464 316230 703520
rect 316454 703464 332422 703520
rect 332646 703464 348706 703520
rect 348930 703464 364898 703520
rect 365122 703464 381090 703520
rect 381314 703464 397374 703520
rect 397598 703464 413566 703520
rect 413790 703464 429758 703520
rect 429982 703464 446042 703520
rect 446266 703464 462234 703520
rect 462458 703464 478426 703520
rect 478650 703464 494710 703520
rect 494934 703464 510902 703520
rect 511126 703464 527094 703520
rect 527318 703464 543378 703520
rect 543602 703464 559570 703520
rect 559794 703464 575762 703520
rect 575986 703464 581422 703520
rect 572 536 581422 703464
rect 710 480 1590 536
rect 1814 480 2786 536
rect 3010 480 3982 536
rect 4206 480 5178 536
rect 5402 480 6374 536
rect 6598 480 7570 536
rect 7794 480 8766 536
rect 8990 480 9962 536
rect 10186 480 11158 536
rect 11382 480 12354 536
rect 12578 480 13550 536
rect 13774 480 14746 536
rect 14970 480 15942 536
rect 16166 480 17138 536
rect 17362 480 18242 536
rect 18466 480 19438 536
rect 19662 480 20634 536
rect 20858 480 21830 536
rect 22054 480 23026 536
rect 23250 480 24222 536
rect 24446 480 25418 536
rect 25642 480 26614 536
rect 26838 480 27810 536
rect 28034 480 29006 536
rect 29230 480 30202 536
rect 30426 480 31398 536
rect 31622 480 32594 536
rect 32818 480 33790 536
rect 34014 480 34894 536
rect 35118 480 36090 536
rect 36314 480 37286 536
rect 37510 480 38482 536
rect 38706 480 39678 536
rect 39902 480 40874 536
rect 41098 480 42070 536
rect 42294 480 43266 536
rect 43490 480 44462 536
rect 44686 480 45658 536
rect 45882 480 46854 536
rect 47078 480 48050 536
rect 48274 480 49246 536
rect 49470 480 50442 536
rect 50666 480 51546 536
rect 51770 480 52742 536
rect 52966 480 53938 536
rect 54162 480 55134 536
rect 55358 480 56330 536
rect 56554 480 57526 536
rect 57750 480 58722 536
rect 58946 480 59918 536
rect 60142 480 61114 536
rect 61338 480 62310 536
rect 62534 480 63506 536
rect 63730 480 64702 536
rect 64926 480 65898 536
rect 66122 480 67094 536
rect 67318 480 68198 536
rect 68422 480 69394 536
rect 69618 480 70590 536
rect 70814 480 71786 536
rect 72010 480 72982 536
rect 73206 480 74178 536
rect 74402 480 75374 536
rect 75598 480 76570 536
rect 76794 480 77766 536
rect 77990 480 78962 536
rect 79186 480 80158 536
rect 80382 480 81354 536
rect 81578 480 82550 536
rect 82774 480 83746 536
rect 83970 480 84850 536
rect 85074 480 86046 536
rect 86270 480 87242 536
rect 87466 480 88438 536
rect 88662 480 89634 536
rect 89858 480 90830 536
rect 91054 480 92026 536
rect 92250 480 93222 536
rect 93446 480 94418 536
rect 94642 480 95614 536
rect 95838 480 96810 536
rect 97034 480 98006 536
rect 98230 480 99202 536
rect 99426 480 100398 536
rect 100622 480 101502 536
rect 101726 480 102698 536
rect 102922 480 103894 536
rect 104118 480 105090 536
rect 105314 480 106286 536
rect 106510 480 107482 536
rect 107706 480 108678 536
rect 108902 480 109874 536
rect 110098 480 111070 536
rect 111294 480 112266 536
rect 112490 480 113462 536
rect 113686 480 114658 536
rect 114882 480 115854 536
rect 116078 480 117050 536
rect 117274 480 118154 536
rect 118378 480 119350 536
rect 119574 480 120546 536
rect 120770 480 121742 536
rect 121966 480 122938 536
rect 123162 480 124134 536
rect 124358 480 125330 536
rect 125554 480 126526 536
rect 126750 480 127722 536
rect 127946 480 128918 536
rect 129142 480 130114 536
rect 130338 480 131310 536
rect 131534 480 132506 536
rect 132730 480 133702 536
rect 133926 480 134806 536
rect 135030 480 136002 536
rect 136226 480 137198 536
rect 137422 480 138394 536
rect 138618 480 139590 536
rect 139814 480 140786 536
rect 141010 480 141982 536
rect 142206 480 143178 536
rect 143402 480 144374 536
rect 144598 480 145570 536
rect 145794 480 146766 536
rect 146990 480 147962 536
rect 148186 480 149158 536
rect 149382 480 150354 536
rect 150578 480 151458 536
rect 151682 480 152654 536
rect 152878 480 153850 536
rect 154074 480 155046 536
rect 155270 480 156242 536
rect 156466 480 157438 536
rect 157662 480 158634 536
rect 158858 480 159830 536
rect 160054 480 161026 536
rect 161250 480 162222 536
rect 162446 480 163418 536
rect 163642 480 164614 536
rect 164838 480 165810 536
rect 166034 480 167006 536
rect 167230 480 168110 536
rect 168334 480 169306 536
rect 169530 480 170502 536
rect 170726 480 171698 536
rect 171922 480 172894 536
rect 173118 480 174090 536
rect 174314 480 175286 536
rect 175510 480 176482 536
rect 176706 480 177678 536
rect 177902 480 178874 536
rect 179098 480 180070 536
rect 180294 480 181266 536
rect 181490 480 182462 536
rect 182686 480 183658 536
rect 183882 480 184762 536
rect 184986 480 185958 536
rect 186182 480 187154 536
rect 187378 480 188350 536
rect 188574 480 189546 536
rect 189770 480 190742 536
rect 190966 480 191938 536
rect 192162 480 193134 536
rect 193358 480 194330 536
rect 194554 480 195526 536
rect 195750 480 196722 536
rect 196946 480 197918 536
rect 198142 480 199114 536
rect 199338 480 200310 536
rect 200534 480 201414 536
rect 201638 480 202610 536
rect 202834 480 203806 536
rect 204030 480 205002 536
rect 205226 480 206198 536
rect 206422 480 207394 536
rect 207618 480 208590 536
rect 208814 480 209786 536
rect 210010 480 210982 536
rect 211206 480 212178 536
rect 212402 480 213374 536
rect 213598 480 214570 536
rect 214794 480 215766 536
rect 215990 480 216962 536
rect 217186 480 218066 536
rect 218290 480 219262 536
rect 219486 480 220458 536
rect 220682 480 221654 536
rect 221878 480 222850 536
rect 223074 480 224046 536
rect 224270 480 225242 536
rect 225466 480 226438 536
rect 226662 480 227634 536
rect 227858 480 228830 536
rect 229054 480 230026 536
rect 230250 480 231222 536
rect 231446 480 232418 536
rect 232642 480 233614 536
rect 233838 480 234718 536
rect 234942 480 235914 536
rect 236138 480 237110 536
rect 237334 480 238306 536
rect 238530 480 239502 536
rect 239726 480 240698 536
rect 240922 480 241894 536
rect 242118 480 243090 536
rect 243314 480 244286 536
rect 244510 480 245482 536
rect 245706 480 246678 536
rect 246902 480 247874 536
rect 248098 480 249070 536
rect 249294 480 250266 536
rect 250490 480 251370 536
rect 251594 480 252566 536
rect 252790 480 253762 536
rect 253986 480 254958 536
rect 255182 480 256154 536
rect 256378 480 257350 536
rect 257574 480 258546 536
rect 258770 480 259742 536
rect 259966 480 260938 536
rect 261162 480 262134 536
rect 262358 480 263330 536
rect 263554 480 264526 536
rect 264750 480 265722 536
rect 265946 480 266918 536
rect 267142 480 268022 536
rect 268246 480 269218 536
rect 269442 480 270414 536
rect 270638 480 271610 536
rect 271834 480 272806 536
rect 273030 480 274002 536
rect 274226 480 275198 536
rect 275422 480 276394 536
rect 276618 480 277590 536
rect 277814 480 278786 536
rect 279010 480 279982 536
rect 280206 480 281178 536
rect 281402 480 282374 536
rect 282598 480 283570 536
rect 283794 480 284674 536
rect 284898 480 285870 536
rect 286094 480 287066 536
rect 287290 480 288262 536
rect 288486 480 289458 536
rect 289682 480 290654 536
rect 290878 480 291850 536
rect 292074 480 293046 536
rect 293270 480 294242 536
rect 294466 480 295438 536
rect 295662 480 296634 536
rect 296858 480 297830 536
rect 298054 480 299026 536
rect 299250 480 300222 536
rect 300446 480 301326 536
rect 301550 480 302522 536
rect 302746 480 303718 536
rect 303942 480 304914 536
rect 305138 480 306110 536
rect 306334 480 307306 536
rect 307530 480 308502 536
rect 308726 480 309698 536
rect 309922 480 310894 536
rect 311118 480 312090 536
rect 312314 480 313286 536
rect 313510 480 314482 536
rect 314706 480 315678 536
rect 315902 480 316874 536
rect 317098 480 317978 536
rect 318202 480 319174 536
rect 319398 480 320370 536
rect 320594 480 321566 536
rect 321790 480 322762 536
rect 322986 480 323958 536
rect 324182 480 325154 536
rect 325378 480 326350 536
rect 326574 480 327546 536
rect 327770 480 328742 536
rect 328966 480 329938 536
rect 330162 480 331134 536
rect 331358 480 332330 536
rect 332554 480 333526 536
rect 333750 480 334630 536
rect 334854 480 335826 536
rect 336050 480 337022 536
rect 337246 480 338218 536
rect 338442 480 339414 536
rect 339638 480 340610 536
rect 340834 480 341806 536
rect 342030 480 343002 536
rect 343226 480 344198 536
rect 344422 480 345394 536
rect 345618 480 346590 536
rect 346814 480 347786 536
rect 348010 480 348982 536
rect 349206 480 350178 536
rect 350402 480 351282 536
rect 351506 480 352478 536
rect 352702 480 353674 536
rect 353898 480 354870 536
rect 355094 480 356066 536
rect 356290 480 357262 536
rect 357486 480 358458 536
rect 358682 480 359654 536
rect 359878 480 360850 536
rect 361074 480 362046 536
rect 362270 480 363242 536
rect 363466 480 364438 536
rect 364662 480 365634 536
rect 365858 480 366830 536
rect 367054 480 367934 536
rect 368158 480 369130 536
rect 369354 480 370326 536
rect 370550 480 371522 536
rect 371746 480 372718 536
rect 372942 480 373914 536
rect 374138 480 375110 536
rect 375334 480 376306 536
rect 376530 480 377502 536
rect 377726 480 378698 536
rect 378922 480 379894 536
rect 380118 480 381090 536
rect 381314 480 382286 536
rect 382510 480 383482 536
rect 383706 480 384586 536
rect 384810 480 385782 536
rect 386006 480 386978 536
rect 387202 480 388174 536
rect 388398 480 389370 536
rect 389594 480 390566 536
rect 390790 480 391762 536
rect 391986 480 392958 536
rect 393182 480 394154 536
rect 394378 480 395350 536
rect 395574 480 396546 536
rect 396770 480 397742 536
rect 397966 480 398938 536
rect 399162 480 400134 536
rect 400358 480 401238 536
rect 401462 480 402434 536
rect 402658 480 403630 536
rect 403854 480 404826 536
rect 405050 480 406022 536
rect 406246 480 407218 536
rect 407442 480 408414 536
rect 408638 480 409610 536
rect 409834 480 410806 536
rect 411030 480 412002 536
rect 412226 480 413198 536
rect 413422 480 414394 536
rect 414618 480 415590 536
rect 415814 480 416786 536
rect 417010 480 417890 536
rect 418114 480 419086 536
rect 419310 480 420282 536
rect 420506 480 421478 536
rect 421702 480 422674 536
rect 422898 480 423870 536
rect 424094 480 425066 536
rect 425290 480 426262 536
rect 426486 480 427458 536
rect 427682 480 428654 536
rect 428878 480 429850 536
rect 430074 480 431046 536
rect 431270 480 432242 536
rect 432466 480 433438 536
rect 433662 480 434542 536
rect 434766 480 435738 536
rect 435962 480 436934 536
rect 437158 480 438130 536
rect 438354 480 439326 536
rect 439550 480 440522 536
rect 440746 480 441718 536
rect 441942 480 442914 536
rect 443138 480 444110 536
rect 444334 480 445306 536
rect 445530 480 446502 536
rect 446726 480 447698 536
rect 447922 480 448894 536
rect 449118 480 450090 536
rect 450314 480 451194 536
rect 451418 480 452390 536
rect 452614 480 453586 536
rect 453810 480 454782 536
rect 455006 480 455978 536
rect 456202 480 457174 536
rect 457398 480 458370 536
rect 458594 480 459566 536
rect 459790 480 460762 536
rect 460986 480 461958 536
rect 462182 480 463154 536
rect 463378 480 464350 536
rect 464574 480 465546 536
rect 465770 480 466742 536
rect 466966 480 467846 536
rect 468070 480 469042 536
rect 469266 480 470238 536
rect 470462 480 471434 536
rect 471658 480 472630 536
rect 472854 480 473826 536
rect 474050 480 475022 536
rect 475246 480 476218 536
rect 476442 480 477414 536
rect 477638 480 478610 536
rect 478834 480 479806 536
rect 480030 480 481002 536
rect 481226 480 482198 536
rect 482422 480 483394 536
rect 483618 480 484498 536
rect 484722 480 485694 536
rect 485918 480 486890 536
rect 487114 480 488086 536
rect 488310 480 489282 536
rect 489506 480 490478 536
rect 490702 480 491674 536
rect 491898 480 492870 536
rect 493094 480 494066 536
rect 494290 480 495262 536
rect 495486 480 496458 536
rect 496682 480 497654 536
rect 497878 480 498850 536
rect 499074 480 500046 536
rect 500270 480 501150 536
rect 501374 480 502346 536
rect 502570 480 503542 536
rect 503766 480 504738 536
rect 504962 480 505934 536
rect 506158 480 507130 536
rect 507354 480 508326 536
rect 508550 480 509522 536
rect 509746 480 510718 536
rect 510942 480 511914 536
rect 512138 480 513110 536
rect 513334 480 514306 536
rect 514530 480 515502 536
rect 515726 480 516698 536
rect 516922 480 517802 536
rect 518026 480 518998 536
rect 519222 480 520194 536
rect 520418 480 521390 536
rect 521614 480 522586 536
rect 522810 480 523782 536
rect 524006 480 524978 536
rect 525202 480 526174 536
rect 526398 480 527370 536
rect 527594 480 528566 536
rect 528790 480 529762 536
rect 529986 480 530958 536
rect 531182 480 532154 536
rect 532378 480 533350 536
rect 533574 480 534454 536
rect 534678 480 535650 536
rect 535874 480 536846 536
rect 537070 480 538042 536
rect 538266 480 539238 536
rect 539462 480 540434 536
rect 540658 480 541630 536
rect 541854 480 542826 536
rect 543050 480 544022 536
rect 544246 480 545218 536
rect 545442 480 546414 536
rect 546638 480 547610 536
rect 547834 480 548806 536
rect 549030 480 550002 536
rect 550226 480 551106 536
rect 551330 480 552302 536
rect 552526 480 553498 536
rect 553722 480 554694 536
rect 554918 480 555890 536
rect 556114 480 557086 536
rect 557310 480 558282 536
rect 558506 480 559478 536
rect 559702 480 560674 536
rect 560898 480 561870 536
rect 562094 480 563066 536
rect 563290 480 564262 536
rect 564486 480 565458 536
rect 565682 480 566654 536
rect 566878 480 567758 536
rect 567982 480 568954 536
rect 569178 480 570150 536
rect 570374 480 571346 536
rect 571570 480 572542 536
rect 572766 480 573738 536
rect 573962 480 574934 536
rect 575158 480 576130 536
rect 576354 480 577326 536
rect 577550 480 578522 536
rect 578746 480 579718 536
rect 579942 480 580914 536
rect 581138 480 581422 536
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 583520 686204 584960 686444
rect -960 682124 480 682364
rect 583520 674508 584960 674748
rect -960 667844 480 668084
rect 583520 662676 584960 662916
rect -960 653428 480 653668
rect 583520 650980 584960 651220
rect -960 639012 480 639252
rect 583520 639284 584960 639524
rect 583520 627588 584960 627828
rect -960 624732 480 624972
rect 583520 615756 584960 615996
rect -960 610316 480 610556
rect 583520 604060 584960 604300
rect -960 595900 480 596140
rect 583520 592364 584960 592604
rect -960 581620 480 581860
rect 583520 580668 584960 580908
rect 583520 568836 584960 569076
rect -960 567204 480 567444
rect 583520 557140 584960 557380
rect -960 552924 480 553164
rect 583520 545444 584960 545684
rect -960 538508 480 538748
rect 583520 533748 584960 533988
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 583520 510220 584960 510460
rect -960 509812 480 510052
rect 583520 498524 584960 498764
rect -960 495396 480 495636
rect 583520 486692 584960 486932
rect -960 480980 480 481220
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 583520 463300 584960 463540
rect -960 452284 480 452524
rect 583520 451604 584960 451844
rect 583520 439772 584960 440012
rect -960 437868 480 438108
rect 583520 428076 584960 428316
rect -960 423588 480 423828
rect 583520 416380 584960 416620
rect -960 409172 480 409412
rect 583520 404684 584960 404924
rect -960 394892 480 395132
rect 583520 392852 584960 393092
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 583520 369460 584960 369700
rect -960 366060 480 366300
rect 583520 357764 584960 358004
rect -960 351780 480 352020
rect 583520 345932 584960 346172
rect -960 337364 480 337604
rect 583520 334236 584960 334476
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 583520 299012 584960 299252
rect -960 294252 480 294492
rect 583520 287316 584960 287556
rect -960 279972 480 280212
rect 583520 275620 584960 275860
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 583520 240396 584960 240636
rect -960 236860 480 237100
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 583520 216868 584960 217108
rect -960 208028 480 208268
rect 583520 205172 584960 205412
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 583520 169948 584960 170188
rect -960 164916 480 165156
rect 583520 158252 584960 158492
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 583520 111332 584960 111572
rect -960 107524 480 107764
rect 583520 99636 584960 99876
rect -960 93108 480 93348
rect 583520 87804 584960 88044
rect -960 78828 480 79068
rect 583520 76108 584960 76348
rect -960 64412 480 64652
rect 583520 64412 584960 64652
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 583520 29188 584960 29428
rect -960 21300 480 21540
rect 583520 17492 584960 17732
rect -960 7020 480 7260
rect 583520 5796 584960 6036
<< obsm3 >>
rect 480 698220 583520 701793
rect 480 697820 583440 698220
rect 480 696860 583520 697820
rect 560 696460 583520 696860
rect 480 686524 583520 696460
rect 480 686124 583440 686524
rect 480 682444 583520 686124
rect 560 682044 583520 682444
rect 480 674828 583520 682044
rect 480 674428 583440 674828
rect 480 668164 583520 674428
rect 560 667764 583520 668164
rect 480 662996 583520 667764
rect 480 662596 583440 662996
rect 480 653748 583520 662596
rect 560 653348 583520 653748
rect 480 651300 583520 653348
rect 480 650900 583440 651300
rect 480 639604 583520 650900
rect 480 639332 583440 639604
rect 560 639204 583440 639332
rect 560 638932 583520 639204
rect 480 627908 583520 638932
rect 480 627508 583440 627908
rect 480 625052 583520 627508
rect 560 624652 583520 625052
rect 480 616076 583520 624652
rect 480 615676 583440 616076
rect 480 610636 583520 615676
rect 560 610236 583520 610636
rect 480 604380 583520 610236
rect 480 603980 583440 604380
rect 480 596220 583520 603980
rect 560 595820 583520 596220
rect 480 592684 583520 595820
rect 480 592284 583440 592684
rect 480 581940 583520 592284
rect 560 581540 583520 581940
rect 480 580988 583520 581540
rect 480 580588 583440 580988
rect 480 569156 583520 580588
rect 480 568756 583440 569156
rect 480 567524 583520 568756
rect 560 567124 583520 567524
rect 480 557460 583520 567124
rect 480 557060 583440 557460
rect 480 553244 583520 557060
rect 560 552844 583520 553244
rect 480 545764 583520 552844
rect 480 545364 583440 545764
rect 480 538828 583520 545364
rect 560 538428 583520 538828
rect 480 534068 583520 538428
rect 480 533668 583440 534068
rect 480 524412 583520 533668
rect 560 524012 583520 524412
rect 480 522236 583520 524012
rect 480 521836 583440 522236
rect 480 510540 583520 521836
rect 480 510140 583440 510540
rect 480 510132 583520 510140
rect 560 509732 583520 510132
rect 480 498844 583520 509732
rect 480 498444 583440 498844
rect 480 495716 583520 498444
rect 560 495316 583520 495716
rect 480 487012 583520 495316
rect 480 486612 583440 487012
rect 480 481300 583520 486612
rect 560 480900 583520 481300
rect 480 475316 583520 480900
rect 480 474916 583440 475316
rect 480 467020 583520 474916
rect 560 466620 583520 467020
rect 480 463620 583520 466620
rect 480 463220 583440 463620
rect 480 452604 583520 463220
rect 560 452204 583520 452604
rect 480 451924 583520 452204
rect 480 451524 583440 451924
rect 480 440092 583520 451524
rect 480 439692 583440 440092
rect 480 438188 583520 439692
rect 560 437788 583520 438188
rect 480 428396 583520 437788
rect 480 427996 583440 428396
rect 480 423908 583520 427996
rect 560 423508 583520 423908
rect 480 416700 583520 423508
rect 480 416300 583440 416700
rect 480 409492 583520 416300
rect 560 409092 583520 409492
rect 480 405004 583520 409092
rect 480 404604 583440 405004
rect 480 395212 583520 404604
rect 560 394812 583520 395212
rect 480 393172 583520 394812
rect 480 392772 583440 393172
rect 480 381476 583520 392772
rect 480 381076 583440 381476
rect 480 380796 583520 381076
rect 560 380396 583520 380796
rect 480 369780 583520 380396
rect 480 369380 583440 369780
rect 480 366380 583520 369380
rect 560 365980 583520 366380
rect 480 358084 583520 365980
rect 480 357684 583440 358084
rect 480 352100 583520 357684
rect 560 351700 583520 352100
rect 480 346252 583520 351700
rect 480 345852 583440 346252
rect 480 337684 583520 345852
rect 560 337284 583520 337684
rect 480 334556 583520 337284
rect 480 334156 583440 334556
rect 480 323268 583520 334156
rect 560 322868 583520 323268
rect 480 322860 583520 322868
rect 480 322460 583440 322860
rect 480 311028 583520 322460
rect 480 310628 583440 311028
rect 480 308988 583520 310628
rect 560 308588 583520 308988
rect 480 299332 583520 308588
rect 480 298932 583440 299332
rect 480 294572 583520 298932
rect 560 294172 583520 294572
rect 480 287636 583520 294172
rect 480 287236 583440 287636
rect 480 280292 583520 287236
rect 560 279892 583520 280292
rect 480 275940 583520 279892
rect 480 275540 583440 275940
rect 480 265876 583520 275540
rect 560 265476 583520 265876
rect 480 264108 583520 265476
rect 480 263708 583440 264108
rect 480 252412 583520 263708
rect 480 252012 583440 252412
rect 480 251460 583520 252012
rect 560 251060 583520 251460
rect 480 240716 583520 251060
rect 480 240316 583440 240716
rect 480 237180 583520 240316
rect 560 236780 583520 237180
rect 480 229020 583520 236780
rect 480 228620 583440 229020
rect 480 222764 583520 228620
rect 560 222364 583520 222764
rect 480 217188 583520 222364
rect 480 216788 583440 217188
rect 480 208348 583520 216788
rect 560 207948 583520 208348
rect 480 205492 583520 207948
rect 480 205092 583440 205492
rect 480 194068 583520 205092
rect 560 193796 583520 194068
rect 560 193668 583440 193796
rect 480 193396 583440 193668
rect 480 182100 583520 193396
rect 480 181700 583440 182100
rect 480 179652 583520 181700
rect 560 179252 583520 179652
rect 480 170268 583520 179252
rect 480 169868 583440 170268
rect 480 165236 583520 169868
rect 560 164836 583520 165236
rect 480 158572 583520 164836
rect 480 158172 583440 158572
rect 480 150956 583520 158172
rect 560 150556 583520 150956
rect 480 146876 583520 150556
rect 480 146476 583440 146876
rect 480 136540 583520 146476
rect 560 136140 583520 136540
rect 480 135044 583520 136140
rect 480 134644 583440 135044
rect 480 123348 583520 134644
rect 480 122948 583440 123348
rect 480 122260 583520 122948
rect 560 121860 583520 122260
rect 480 111652 583520 121860
rect 480 111252 583440 111652
rect 480 107844 583520 111252
rect 560 107444 583520 107844
rect 480 99956 583520 107444
rect 480 99556 583440 99956
rect 480 93428 583520 99556
rect 560 93028 583520 93428
rect 480 88124 583520 93028
rect 480 87724 583440 88124
rect 480 79148 583520 87724
rect 560 78748 583520 79148
rect 480 76428 583520 78748
rect 480 76028 583440 76428
rect 480 64732 583520 76028
rect 560 64332 583440 64732
rect 480 53036 583520 64332
rect 480 52636 583440 53036
rect 480 50316 583520 52636
rect 560 49916 583520 50316
rect 480 41204 583520 49916
rect 480 40804 583440 41204
rect 480 36036 583520 40804
rect 560 35636 583520 36036
rect 480 29508 583520 35636
rect 480 29108 583440 29508
rect 480 21620 583520 29108
rect 560 21220 583520 21620
rect 480 17812 583520 21220
rect 480 17412 583440 17812
rect 480 7340 583520 17412
rect 560 6940 583520 7340
rect 480 6116 583520 6940
rect 480 5716 583440 6116
rect 480 2143 583520 5716
<< metal4 >>
rect -8576 -7504 -7976 711440
rect -7636 -6564 -7036 710500
rect -6696 -5624 -6096 709560
rect -5756 -4684 -5156 708620
rect -4816 -3744 -4216 707680
rect -3876 -2804 -3276 706740
rect -2936 -1864 -2336 705800
rect -1996 -924 -1396 704860
rect 804 -1864 1404 705800
rect 4404 693500 5004 707680
rect 8004 693500 8604 709560
rect 11604 693500 12204 711440
rect 18804 693452 19404 705800
rect 22404 693500 23004 707680
rect 26004 693500 26604 709560
rect 29604 693500 30204 711440
rect 36804 693452 37404 705800
rect 40404 693500 41004 707680
rect 44004 693500 44604 709560
rect 47604 693500 48204 711440
rect 54804 693452 55404 705800
rect 58404 693500 59004 707680
rect 62004 693500 62604 709560
rect 65604 693500 66204 711440
rect 72804 693452 73404 705800
rect 76404 693500 77004 707680
rect 80004 693500 80604 709560
rect 83604 693500 84204 711440
rect 90804 693452 91404 705800
rect 94404 693500 95004 707680
rect 98004 693500 98604 709560
rect 101604 693500 102204 711440
rect 108804 693452 109404 705800
rect 112404 693500 113004 707680
rect 116004 693500 116604 709560
rect 119604 693500 120204 711440
rect 126804 693452 127404 705800
rect 130404 693500 131004 707680
rect 134004 693500 134604 709560
rect 137604 693500 138204 711440
rect 144804 693452 145404 705800
rect 148404 693500 149004 707680
rect 152004 693500 152604 709560
rect 155604 693500 156204 711440
rect 162804 693452 163404 705800
rect 166404 693500 167004 707680
rect 170004 693500 170604 709560
rect 173604 693500 174204 711440
rect 180804 693452 181404 705800
rect 184404 693500 185004 707680
rect 188004 693500 188604 709560
rect 191604 693500 192204 711440
rect 198804 693452 199404 705800
rect 202404 693500 203004 707680
rect 206004 693500 206604 709560
rect 209604 693500 210204 711440
rect 216804 693452 217404 705800
rect 220404 693500 221004 707680
rect 224004 693500 224604 709560
rect 227604 693500 228204 711440
rect 234804 693452 235404 705800
rect 238404 693500 239004 707680
rect 242004 693500 242604 709560
rect 245604 693500 246204 711440
rect 252804 693452 253404 705800
rect 256404 693500 257004 707680
rect 260004 693500 260604 709560
rect 263604 693500 264204 711440
rect 270804 693452 271404 705800
rect 274404 693500 275004 707680
rect 278004 693500 278604 709560
rect 281604 693500 282204 711440
rect 288804 693452 289404 705800
rect 292404 693500 293004 707680
rect 296004 693500 296604 709560
rect 299604 693500 300204 711440
rect 306804 693452 307404 705800
rect 310404 693500 311004 707680
rect 314004 693500 314604 709560
rect 317604 693500 318204 711440
rect 324804 693452 325404 705800
rect 328404 693500 329004 707680
rect 332004 693500 332604 709560
rect 335604 693500 336204 711440
rect 342804 693452 343404 705800
rect 346404 693500 347004 707680
rect 350004 693500 350604 709560
rect 353604 693500 354204 711440
rect 360804 693452 361404 705800
rect 364404 693500 365004 707680
rect 368004 693500 368604 709560
rect 371604 693500 372204 711440
rect 378804 693452 379404 705800
rect 382404 693500 383004 707680
rect 386004 693500 386604 709560
rect 389604 693500 390204 711440
rect 396804 693452 397404 705800
rect 400404 693500 401004 707680
rect 404004 693500 404604 709560
rect 407604 693500 408204 711440
rect 414804 693452 415404 705800
rect 418404 693500 419004 707680
rect 422004 693500 422604 709560
rect 425604 693500 426204 711440
rect 432804 693452 433404 705800
rect 436404 693500 437004 707680
rect 440004 693500 440604 709560
rect 443604 693500 444204 711440
rect 450804 693452 451404 705800
rect 454404 693500 455004 707680
rect 458004 693500 458604 709560
rect 461604 693500 462204 711440
rect 468804 693452 469404 705800
rect 472404 693500 473004 707680
rect 476004 693500 476604 709560
rect 479604 693500 480204 711440
rect 486804 693452 487404 705800
rect 490404 693500 491004 707680
rect 494004 693500 494604 709560
rect 497604 693500 498204 711440
rect 504804 693452 505404 705800
rect 508404 693500 509004 707680
rect 512004 693500 512604 709560
rect 515604 693500 516204 711440
rect 522804 693452 523404 705800
rect 526404 693500 527004 707680
rect 530004 693500 530604 709560
rect 533604 693500 534204 711440
rect 540804 693452 541404 705800
rect 544404 693500 545004 707680
rect 548004 693500 548604 709560
rect 551604 693500 552204 711440
rect 558804 693452 559404 705800
rect 562404 693500 563004 707680
rect 566004 693500 566604 709560
rect 569604 693500 570204 711440
rect 576804 693452 577404 705800
rect 580404 693500 581004 707680
rect 4404 493500 5004 534500
rect 8004 493500 8604 534500
rect 11604 493500 12204 534500
rect 18804 493452 19404 534548
rect 22404 493500 23004 534500
rect 26004 493500 26604 534500
rect 29604 493500 30204 534500
rect 36804 493452 37404 534548
rect 40404 493500 41004 534500
rect 44004 493500 44604 534500
rect 47604 493500 48204 534500
rect 54804 493452 55404 534548
rect 58404 493500 59004 534500
rect 62004 493500 62604 534500
rect 65604 493500 66204 534500
rect 72804 493452 73404 534548
rect 76404 493500 77004 534500
rect 80004 493500 80604 534500
rect 83604 493500 84204 534500
rect 90804 493452 91404 534548
rect 94404 493500 95004 534500
rect 98004 493500 98604 534500
rect 101604 493500 102204 534500
rect 108804 493452 109404 534548
rect 112404 493500 113004 534500
rect 116004 493500 116604 534500
rect 119604 493500 120204 534500
rect 126804 493452 127404 534548
rect 130404 493500 131004 534500
rect 134004 493500 134604 534500
rect 137604 493500 138204 534500
rect 144804 493452 145404 534548
rect 148404 493500 149004 534500
rect 152004 493500 152604 534500
rect 155604 493500 156204 534500
rect 4404 249500 5004 338500
rect 8004 249500 8604 338500
rect 11604 249500 12204 338500
rect 18804 249452 19404 338548
rect 22404 249500 23004 338500
rect 26004 249500 26604 338500
rect 29604 249500 30204 338500
rect 36804 249452 37404 338548
rect 40404 249500 41004 338500
rect 44004 249500 44604 338500
rect 47604 249500 48204 338500
rect 54804 249452 55404 338548
rect 58404 249500 59004 338500
rect 62004 249500 62604 338500
rect 65604 249500 66204 338500
rect 72804 249452 73404 338548
rect 76404 249500 77004 338500
rect 80004 249500 80604 338500
rect 83604 249500 84204 338500
rect 90804 249452 91404 338548
rect 94404 249500 95004 338500
rect 98004 249500 98604 338500
rect 101604 249500 102204 338500
rect 108804 249452 109404 338548
rect 112404 249500 113004 338500
rect 116004 249500 116604 338500
rect 119604 249500 120204 338500
rect 126804 249452 127404 338548
rect 130404 249500 131004 338500
rect 134004 249500 134604 338500
rect 137604 249500 138204 338500
rect 144804 249452 145404 338548
rect 148404 249500 149004 338500
rect 152004 249500 152604 338500
rect 155604 249500 156204 338500
rect 162804 249452 163404 534548
rect 166404 249500 167004 534500
rect 170004 249500 170604 534500
rect 173604 249500 174204 534500
rect 180804 249452 181404 534548
rect 184404 249500 185004 534500
rect 188004 249500 188604 534500
rect 191604 249500 192204 534500
rect 198804 249452 199404 534548
rect 202404 249500 203004 534500
rect 206004 249500 206604 534500
rect 209604 249500 210204 534500
rect 216804 249452 217404 534548
rect 220404 249500 221004 534500
rect 224004 249500 224604 534500
rect 227604 249500 228204 534500
rect 234804 249452 235404 534548
rect 238404 249500 239004 534500
rect 4404 -3744 5004 10500
rect 8004 -5624 8604 10500
rect 11604 -7504 12204 10500
rect 18804 -1864 19404 10548
rect 22404 -3744 23004 10500
rect 26004 -5624 26604 10500
rect 29604 -7504 30204 10500
rect 36804 -1864 37404 10548
rect 40404 -3744 41004 10500
rect 44004 -5624 44604 10500
rect 47604 -7504 48204 10500
rect 54804 -1864 55404 10548
rect 58404 -3744 59004 10500
rect 62004 -5624 62604 10500
rect 65604 -7504 66204 10500
rect 72804 -1864 73404 10548
rect 76404 -3744 77004 10500
rect 80004 -5624 80604 10500
rect 83604 -7504 84204 10500
rect 90804 -1864 91404 10548
rect 94404 -3744 95004 10500
rect 98004 -5624 98604 10500
rect 101604 -7504 102204 10500
rect 108804 -1864 109404 10548
rect 112404 -3744 113004 10500
rect 116004 -5624 116604 10500
rect 119604 -7504 120204 10500
rect 126804 -1864 127404 10548
rect 130404 -3744 131004 10500
rect 134004 -5624 134604 10500
rect 137604 -7504 138204 10500
rect 144804 -1864 145404 10548
rect 148404 -3744 149004 10500
rect 152004 -5624 152604 10500
rect 155604 -7504 156204 10500
rect 162804 -1864 163404 10548
rect 166404 -3744 167004 10500
rect 170004 -5624 170604 10500
rect 173604 -7504 174204 10500
rect 180804 -1864 181404 10548
rect 184404 -3744 185004 10500
rect 188004 -5624 188604 10500
rect 191604 -7504 192204 10500
rect 198804 -1864 199404 10548
rect 202404 -3744 203004 10500
rect 206004 -5624 206604 10500
rect 209604 -7504 210204 10500
rect 216804 -1864 217404 10548
rect 220404 -3744 221004 10500
rect 224004 -5624 224604 10500
rect 227604 -7504 228204 10500
rect 234804 -1864 235404 10548
rect 238404 -3744 239004 10500
rect 242004 -5624 242604 534500
rect 245604 -7504 246204 534500
rect 252804 -1864 253404 534548
rect 256404 -3744 257004 534500
rect 260004 -5624 260604 534500
rect 263604 -7504 264204 534500
rect 270804 -1864 271404 534548
rect 274404 -3744 275004 534500
rect 278004 -5624 278604 534500
rect 281604 -7504 282204 534500
rect 288804 -1864 289404 534548
rect 292404 -3744 293004 534500
rect 296004 -5624 296604 534500
rect 299604 -7504 300204 534500
rect 306804 -1864 307404 534548
rect 310404 -3744 311004 534500
rect 314004 -5624 314604 534500
rect 317604 -7504 318204 534500
rect 324804 -1864 325404 534548
rect 328404 -3744 329004 534500
rect 332004 -5624 332604 534500
rect 335604 -7504 336204 534500
rect 342804 249452 343404 534548
rect 346404 249500 347004 534500
rect 350004 249500 350604 534500
rect 353604 249500 354204 534500
rect 360804 249452 361404 534548
rect 364404 249500 365004 534500
rect 368004 249500 368604 534500
rect 371604 249500 372204 534500
rect 378804 249452 379404 534548
rect 382404 249500 383004 534500
rect 386004 249500 386604 534500
rect 389604 249500 390204 534500
rect 396804 249452 397404 534548
rect 400404 249500 401004 534500
rect 404004 249500 404604 534500
rect 407604 249500 408204 534500
rect 414804 503452 415404 534548
rect 418404 503500 419004 534500
rect 422004 503500 422604 534500
rect 425604 503500 426204 534500
rect 432804 503452 433404 534548
rect 436404 503500 437004 534500
rect 440004 503500 440604 534500
rect 443604 503500 444204 534500
rect 450804 503452 451404 534548
rect 454404 503500 455004 534500
rect 458004 503500 458604 534500
rect 461604 503500 462204 534500
rect 468804 503452 469404 534548
rect 472404 503500 473004 534500
rect 476004 503500 476604 534500
rect 479604 503500 480204 534500
rect 486804 503452 487404 534548
rect 490404 503500 491004 534500
rect 494004 503500 494604 534500
rect 497604 503500 498204 534500
rect 504804 503452 505404 534548
rect 508404 503500 509004 534500
rect 512004 503500 512604 534500
rect 515604 503500 516204 534500
rect 522804 503452 523404 534548
rect 526404 503500 527004 534500
rect 530004 503500 530604 534500
rect 533604 503500 534204 534500
rect 540804 503452 541404 534548
rect 544404 503500 545004 534500
rect 548004 503500 548604 534500
rect 551604 503500 552204 534500
rect 558804 503452 559404 534548
rect 562404 503500 563004 534500
rect 566004 503500 566604 534500
rect 569604 503500 570204 534500
rect 576804 503452 577404 534548
rect 580404 503500 581004 534500
rect 414804 249452 415404 334548
rect 418404 249500 419004 334500
rect 422004 249500 422604 334500
rect 425604 249500 426204 334500
rect 432804 249452 433404 334548
rect 436404 249500 437004 334500
rect 440004 249500 440604 334500
rect 443604 249500 444204 334500
rect 450804 249452 451404 334548
rect 454404 249500 455004 334500
rect 458004 249500 458604 334500
rect 461604 249500 462204 334500
rect 468804 249452 469404 334548
rect 472404 249500 473004 334500
rect 476004 249500 476604 334500
rect 479604 249500 480204 334500
rect 486804 249452 487404 334548
rect 490404 249500 491004 334500
rect 494004 249500 494604 334500
rect 497604 249500 498204 334500
rect 504804 249452 505404 334548
rect 508404 249500 509004 334500
rect 512004 249500 512604 334500
rect 515604 249500 516204 334500
rect 522804 249452 523404 334548
rect 526404 249500 527004 334500
rect 530004 249500 530604 334500
rect 533604 249500 534204 334500
rect 540804 249452 541404 334548
rect 544404 249500 545004 334500
rect 548004 249500 548604 334500
rect 551604 249500 552204 334500
rect 558804 249452 559404 334548
rect 562404 249500 563004 334500
rect 566004 249500 566604 334500
rect 569604 249500 570204 334500
rect 576804 249452 577404 334548
rect 580404 249500 581004 334500
rect 342804 -1864 343404 10548
rect 346404 -3744 347004 10500
rect 350004 -5624 350604 10500
rect 353604 -7504 354204 10500
rect 360804 -1864 361404 10548
rect 364404 -3744 365004 10500
rect 368004 -5624 368604 10500
rect 371604 -7504 372204 10500
rect 378804 -1864 379404 10548
rect 382404 -3744 383004 10500
rect 386004 -5624 386604 10500
rect 389604 -7504 390204 10500
rect 396804 -1864 397404 10548
rect 400404 -3744 401004 10500
rect 404004 -5624 404604 10500
rect 407604 -7504 408204 10500
rect 414804 -1864 415404 10548
rect 418404 -3744 419004 10500
rect 422004 -5624 422604 10500
rect 425604 -7504 426204 10500
rect 432804 -1864 433404 10548
rect 436404 -3744 437004 10500
rect 440004 -5624 440604 10500
rect 443604 -7504 444204 10500
rect 450804 -1864 451404 10548
rect 454404 -3744 455004 10500
rect 458004 -5624 458604 10500
rect 461604 -7504 462204 10500
rect 468804 -1864 469404 10548
rect 472404 -3744 473004 10500
rect 476004 -5624 476604 10500
rect 479604 -7504 480204 10500
rect 486804 -1864 487404 10548
rect 490404 -3744 491004 10500
rect 494004 -5624 494604 10500
rect 497604 -7504 498204 10500
rect 504804 -1864 505404 10548
rect 508404 -3744 509004 10500
rect 512004 -5624 512604 10500
rect 515604 -7504 516204 10500
rect 522804 -1864 523404 10548
rect 526404 -3744 527004 10500
rect 530004 -5624 530604 10500
rect 533604 -7504 534204 10500
rect 540804 -1864 541404 10548
rect 544404 -3744 545004 10500
rect 548004 -5624 548604 10500
rect 551604 -7504 552204 10500
rect 558804 -1864 559404 10548
rect 562404 -3744 563004 10500
rect 566004 -5624 566604 10500
rect 569604 -7504 570204 10500
rect 576804 -1864 577404 10548
rect 580404 -3744 581004 10500
rect 585320 -924 585920 704860
rect 586260 -1864 586860 705800
rect 587200 -2804 587800 706740
rect 588140 -3744 588740 707680
rect 589080 -4684 589680 708620
rect 590020 -5624 590620 709560
rect 590960 -6564 591560 710500
rect 591900 -7504 592500 711440
<< obsm4 >>
rect 15555 534628 569797 681680
rect 15555 493372 18724 534628
rect 19484 534580 36724 534628
rect 19484 493420 22324 534580
rect 23084 493420 25924 534580
rect 26684 493420 29524 534580
rect 30284 493420 36724 534580
rect 37484 534580 54724 534628
rect 19484 493372 36724 493420
rect 37484 493420 40324 534580
rect 41084 493420 43924 534580
rect 44684 493420 47524 534580
rect 48284 493420 54724 534580
rect 55484 534580 72724 534628
rect 37484 493372 54724 493420
rect 55484 493420 58324 534580
rect 59084 493420 61924 534580
rect 62684 493420 65524 534580
rect 66284 493420 72724 534580
rect 73484 534580 90724 534628
rect 55484 493372 72724 493420
rect 73484 493420 76324 534580
rect 77084 493420 79924 534580
rect 80684 493420 83524 534580
rect 84284 493420 90724 534580
rect 91484 534580 108724 534628
rect 73484 493372 90724 493420
rect 91484 493420 94324 534580
rect 95084 493420 97924 534580
rect 98684 493420 101524 534580
rect 102284 493420 108724 534580
rect 109484 534580 126724 534628
rect 91484 493372 108724 493420
rect 109484 493420 112324 534580
rect 113084 493420 115924 534580
rect 116684 493420 119524 534580
rect 120284 493420 126724 534580
rect 127484 534580 144724 534628
rect 109484 493372 126724 493420
rect 127484 493420 130324 534580
rect 131084 493420 133924 534580
rect 134684 493420 137524 534580
rect 138284 493420 144724 534580
rect 145484 534580 162724 534628
rect 127484 493372 144724 493420
rect 145484 493420 148324 534580
rect 149084 493420 151924 534580
rect 152684 493420 155524 534580
rect 156284 493420 162724 534580
rect 163484 534580 180724 534628
rect 145484 493372 162724 493420
rect 15555 338628 162724 493372
rect 15555 249372 18724 338628
rect 19484 338580 36724 338628
rect 19484 249420 22324 338580
rect 23084 249420 25924 338580
rect 26684 249420 29524 338580
rect 30284 249420 36724 338580
rect 37484 338580 54724 338628
rect 19484 249372 36724 249420
rect 37484 249420 40324 338580
rect 41084 249420 43924 338580
rect 44684 249420 47524 338580
rect 48284 249420 54724 338580
rect 55484 338580 72724 338628
rect 37484 249372 54724 249420
rect 55484 249420 58324 338580
rect 59084 249420 61924 338580
rect 62684 249420 65524 338580
rect 66284 249420 72724 338580
rect 73484 338580 90724 338628
rect 55484 249372 72724 249420
rect 73484 249420 76324 338580
rect 77084 249420 79924 338580
rect 80684 249420 83524 338580
rect 84284 249420 90724 338580
rect 91484 338580 108724 338628
rect 73484 249372 90724 249420
rect 91484 249420 94324 338580
rect 95084 249420 97924 338580
rect 98684 249420 101524 338580
rect 102284 249420 108724 338580
rect 109484 338580 126724 338628
rect 91484 249372 108724 249420
rect 109484 249420 112324 338580
rect 113084 249420 115924 338580
rect 116684 249420 119524 338580
rect 120284 249420 126724 338580
rect 127484 338580 144724 338628
rect 109484 249372 126724 249420
rect 127484 249420 130324 338580
rect 131084 249420 133924 338580
rect 134684 249420 137524 338580
rect 138284 249420 144724 338580
rect 145484 338580 162724 338628
rect 127484 249372 144724 249420
rect 145484 249420 148324 338580
rect 149084 249420 151924 338580
rect 152684 249420 155524 338580
rect 156284 249420 162724 338580
rect 145484 249372 162724 249420
rect 163484 249420 166324 534580
rect 167084 249420 169924 534580
rect 170684 249420 173524 534580
rect 174284 249420 180724 534580
rect 181484 534580 198724 534628
rect 163484 249372 180724 249420
rect 181484 249420 184324 534580
rect 185084 249420 187924 534580
rect 188684 249420 191524 534580
rect 192284 249420 198724 534580
rect 199484 534580 216724 534628
rect 181484 249372 198724 249420
rect 199484 249420 202324 534580
rect 203084 249420 205924 534580
rect 206684 249420 209524 534580
rect 210284 249420 216724 534580
rect 217484 534580 234724 534628
rect 199484 249372 216724 249420
rect 217484 249420 220324 534580
rect 221084 249420 223924 534580
rect 224684 249420 227524 534580
rect 228284 249420 234724 534580
rect 235484 534580 252724 534628
rect 217484 249372 234724 249420
rect 235484 249420 238324 534580
rect 239084 249420 241924 534580
rect 235484 249372 241924 249420
rect 15555 10628 241924 249372
rect 15555 3299 18724 10628
rect 19484 10580 36724 10628
rect 19484 3299 22324 10580
rect 23084 3299 25924 10580
rect 26684 3299 29524 10580
rect 30284 3299 36724 10580
rect 37484 10580 54724 10628
rect 37484 3299 40324 10580
rect 41084 3299 43924 10580
rect 44684 3299 47524 10580
rect 48284 3299 54724 10580
rect 55484 10580 72724 10628
rect 55484 3299 58324 10580
rect 59084 3299 61924 10580
rect 62684 3299 65524 10580
rect 66284 3299 72724 10580
rect 73484 10580 90724 10628
rect 73484 3299 76324 10580
rect 77084 3299 79924 10580
rect 80684 3299 83524 10580
rect 84284 3299 90724 10580
rect 91484 10580 108724 10628
rect 91484 3299 94324 10580
rect 95084 3299 97924 10580
rect 98684 3299 101524 10580
rect 102284 3299 108724 10580
rect 109484 10580 126724 10628
rect 109484 3299 112324 10580
rect 113084 3299 115924 10580
rect 116684 3299 119524 10580
rect 120284 3299 126724 10580
rect 127484 10580 144724 10628
rect 127484 3299 130324 10580
rect 131084 3299 133924 10580
rect 134684 3299 137524 10580
rect 138284 3299 144724 10580
rect 145484 10580 162724 10628
rect 145484 3299 148324 10580
rect 149084 3299 151924 10580
rect 152684 3299 155524 10580
rect 156284 3299 162724 10580
rect 163484 10580 180724 10628
rect 163484 3299 166324 10580
rect 167084 3299 169924 10580
rect 170684 3299 173524 10580
rect 174284 3299 180724 10580
rect 181484 10580 198724 10628
rect 181484 3299 184324 10580
rect 185084 3299 187924 10580
rect 188684 3299 191524 10580
rect 192284 3299 198724 10580
rect 199484 10580 216724 10628
rect 199484 3299 202324 10580
rect 203084 3299 205924 10580
rect 206684 3299 209524 10580
rect 210284 3299 216724 10580
rect 217484 10580 234724 10628
rect 217484 3299 220324 10580
rect 221084 3299 223924 10580
rect 224684 3299 227524 10580
rect 228284 3299 234724 10580
rect 235484 10580 241924 10628
rect 235484 3299 238324 10580
rect 239084 3299 241924 10580
rect 242684 3299 245524 534580
rect 246284 3299 252724 534580
rect 253484 534580 270724 534628
rect 253484 3299 256324 534580
rect 257084 3299 259924 534580
rect 260684 3299 263524 534580
rect 264284 3299 270724 534580
rect 271484 534580 288724 534628
rect 271484 3299 274324 534580
rect 275084 3299 277924 534580
rect 278684 3299 281524 534580
rect 282284 3299 288724 534580
rect 289484 534580 306724 534628
rect 289484 3299 292324 534580
rect 293084 3299 295924 534580
rect 296684 3299 299524 534580
rect 300284 3299 306724 534580
rect 307484 534580 324724 534628
rect 307484 3299 310324 534580
rect 311084 3299 313924 534580
rect 314684 3299 317524 534580
rect 318284 3299 324724 534580
rect 325484 534580 342724 534628
rect 325484 3299 328324 534580
rect 329084 3299 331924 534580
rect 332684 3299 335524 534580
rect 336284 249372 342724 534580
rect 343484 534580 360724 534628
rect 343484 249420 346324 534580
rect 347084 249420 349924 534580
rect 350684 249420 353524 534580
rect 354284 249420 360724 534580
rect 361484 534580 378724 534628
rect 343484 249372 360724 249420
rect 361484 249420 364324 534580
rect 365084 249420 367924 534580
rect 368684 249420 371524 534580
rect 372284 249420 378724 534580
rect 379484 534580 396724 534628
rect 361484 249372 378724 249420
rect 379484 249420 382324 534580
rect 383084 249420 385924 534580
rect 386684 249420 389524 534580
rect 390284 249420 396724 534580
rect 397484 534580 414724 534628
rect 379484 249372 396724 249420
rect 397484 249420 400324 534580
rect 401084 249420 403924 534580
rect 404684 249420 407524 534580
rect 408284 503372 414724 534580
rect 415484 534580 432724 534628
rect 415484 503420 418324 534580
rect 419084 503420 421924 534580
rect 422684 503420 425524 534580
rect 426284 503420 432724 534580
rect 433484 534580 450724 534628
rect 415484 503372 432724 503420
rect 433484 503420 436324 534580
rect 437084 503420 439924 534580
rect 440684 503420 443524 534580
rect 444284 503420 450724 534580
rect 451484 534580 468724 534628
rect 433484 503372 450724 503420
rect 451484 503420 454324 534580
rect 455084 503420 457924 534580
rect 458684 503420 461524 534580
rect 462284 503420 468724 534580
rect 469484 534580 486724 534628
rect 451484 503372 468724 503420
rect 469484 503420 472324 534580
rect 473084 503420 475924 534580
rect 476684 503420 479524 534580
rect 480284 503420 486724 534580
rect 487484 534580 504724 534628
rect 469484 503372 486724 503420
rect 487484 503420 490324 534580
rect 491084 503420 493924 534580
rect 494684 503420 497524 534580
rect 498284 503420 504724 534580
rect 505484 534580 522724 534628
rect 487484 503372 504724 503420
rect 505484 503420 508324 534580
rect 509084 503420 511924 534580
rect 512684 503420 515524 534580
rect 516284 503420 522724 534580
rect 523484 534580 540724 534628
rect 505484 503372 522724 503420
rect 523484 503420 526324 534580
rect 527084 503420 529924 534580
rect 530684 503420 533524 534580
rect 534284 503420 540724 534580
rect 541484 534580 558724 534628
rect 523484 503372 540724 503420
rect 541484 503420 544324 534580
rect 545084 503420 547924 534580
rect 548684 503420 551524 534580
rect 552284 503420 558724 534580
rect 559484 534580 569797 534628
rect 541484 503372 558724 503420
rect 559484 503420 562324 534580
rect 563084 503420 565924 534580
rect 566684 503420 569524 534580
rect 559484 503372 569797 503420
rect 408284 334628 569797 503372
rect 408284 249420 414724 334628
rect 415484 334580 432724 334628
rect 397484 249372 414724 249420
rect 415484 249420 418324 334580
rect 419084 249420 421924 334580
rect 422684 249420 425524 334580
rect 426284 249420 432724 334580
rect 433484 334580 450724 334628
rect 415484 249372 432724 249420
rect 433484 249420 436324 334580
rect 437084 249420 439924 334580
rect 440684 249420 443524 334580
rect 444284 249420 450724 334580
rect 451484 334580 468724 334628
rect 433484 249372 450724 249420
rect 451484 249420 454324 334580
rect 455084 249420 457924 334580
rect 458684 249420 461524 334580
rect 462284 249420 468724 334580
rect 469484 334580 486724 334628
rect 451484 249372 468724 249420
rect 469484 249420 472324 334580
rect 473084 249420 475924 334580
rect 476684 249420 479524 334580
rect 480284 249420 486724 334580
rect 487484 334580 504724 334628
rect 469484 249372 486724 249420
rect 487484 249420 490324 334580
rect 491084 249420 493924 334580
rect 494684 249420 497524 334580
rect 498284 249420 504724 334580
rect 505484 334580 522724 334628
rect 487484 249372 504724 249420
rect 505484 249420 508324 334580
rect 509084 249420 511924 334580
rect 512684 249420 515524 334580
rect 516284 249420 522724 334580
rect 523484 334580 540724 334628
rect 505484 249372 522724 249420
rect 523484 249420 526324 334580
rect 527084 249420 529924 334580
rect 530684 249420 533524 334580
rect 534284 249420 540724 334580
rect 541484 334580 558724 334628
rect 523484 249372 540724 249420
rect 541484 249420 544324 334580
rect 545084 249420 547924 334580
rect 548684 249420 551524 334580
rect 552284 249420 558724 334580
rect 559484 334580 569797 334628
rect 541484 249372 558724 249420
rect 559484 249420 562324 334580
rect 563084 249420 565924 334580
rect 566684 249420 569524 334580
rect 559484 249372 569797 249420
rect 336284 10628 569797 249372
rect 336284 3299 342724 10628
rect 343484 10580 360724 10628
rect 343484 3299 346324 10580
rect 347084 3299 349924 10580
rect 350684 3299 353524 10580
rect 354284 3299 360724 10580
rect 361484 10580 378724 10628
rect 361484 3299 364324 10580
rect 365084 3299 367924 10580
rect 368684 3299 371524 10580
rect 372284 3299 378724 10580
rect 379484 10580 396724 10628
rect 379484 3299 382324 10580
rect 383084 3299 385924 10580
rect 386684 3299 389524 10580
rect 390284 3299 396724 10580
rect 397484 10580 414724 10628
rect 397484 3299 400324 10580
rect 401084 3299 403924 10580
rect 404684 3299 407524 10580
rect 408284 3299 414724 10580
rect 415484 10580 432724 10628
rect 415484 3299 418324 10580
rect 419084 3299 421924 10580
rect 422684 3299 425524 10580
rect 426284 3299 432724 10580
rect 433484 10580 450724 10628
rect 433484 3299 436324 10580
rect 437084 3299 439924 10580
rect 440684 3299 443524 10580
rect 444284 3299 450724 10580
rect 451484 10580 468724 10628
rect 451484 3299 454324 10580
rect 455084 3299 457924 10580
rect 458684 3299 461524 10580
rect 462284 3299 468724 10580
rect 469484 10580 486724 10628
rect 469484 3299 472324 10580
rect 473084 3299 475924 10580
rect 476684 3299 479524 10580
rect 480284 3299 486724 10580
rect 487484 10580 504724 10628
rect 487484 3299 490324 10580
rect 491084 3299 493924 10580
rect 494684 3299 497524 10580
rect 498284 3299 504724 10580
rect 505484 10580 522724 10628
rect 505484 3299 508324 10580
rect 509084 3299 511924 10580
rect 512684 3299 515524 10580
rect 516284 3299 522724 10580
rect 523484 10580 540724 10628
rect 523484 3299 526324 10580
rect 527084 3299 529924 10580
rect 530684 3299 533524 10580
rect 534284 3299 540724 10580
rect 541484 10580 558724 10628
rect 541484 3299 544324 10580
rect 545084 3299 547924 10580
rect 548684 3299 551524 10580
rect 552284 3299 558724 10580
rect 559484 10580 569797 10628
rect 559484 3299 562324 10580
rect 563084 3299 565924 10580
rect 566684 3299 569524 10580
<< metal5 >>
rect -8576 710840 592500 711440
rect -7636 709900 591560 710500
rect -6696 708960 590620 709560
rect -5756 708020 589680 708620
rect -4816 707080 588740 707680
rect -3876 706140 587800 706740
rect -2936 705200 586860 705800
rect -1996 704260 585920 704860
rect -8576 696676 592500 697276
rect -6696 693076 590620 693676
rect -4816 689476 588740 690076
rect -2936 685828 586860 686428
rect -8576 678676 592500 679276
rect -6696 675076 590620 675676
rect -4816 671476 588740 672076
rect -2936 667828 586860 668428
rect -8576 660676 592500 661276
rect -6696 657076 590620 657676
rect -4816 653476 588740 654076
rect -2936 649828 586860 650428
rect -8576 642676 592500 643276
rect -6696 639076 590620 639676
rect -4816 635476 588740 636076
rect -2936 631828 586860 632428
rect -8576 624676 592500 625276
rect -6696 621076 590620 621676
rect -4816 617476 588740 618076
rect -2936 613828 586860 614428
rect -8576 606676 592500 607276
rect -6696 603076 590620 603676
rect -4816 599476 588740 600076
rect -2936 595828 586860 596428
rect -8576 588676 592500 589276
rect -6696 585076 590620 585676
rect -4816 581476 588740 582076
rect -2936 577828 586860 578428
rect -8576 570676 592500 571276
rect -6696 567076 590620 567676
rect -4816 563476 588740 564076
rect -2936 559828 586860 560428
rect -8576 552676 592500 553276
rect -6696 549076 590620 549676
rect -4816 545476 588740 546076
rect -2936 541828 586860 542428
rect -8576 534676 592500 535276
rect -6696 531076 590620 531676
rect -4816 527476 588740 528076
rect -2936 523828 586860 524428
rect -8576 516676 592500 517276
rect -6696 513076 590620 513676
rect -4816 509476 588740 510076
rect -2936 505828 586860 506428
rect -8576 498676 592500 499276
rect -6696 495076 590620 495676
rect -4816 491476 588740 492076
rect -2936 487828 586860 488428
rect -8576 480676 592500 481276
rect -6696 477076 590620 477676
rect -4816 473476 588740 474076
rect -2936 469828 586860 470428
rect -8576 462676 592500 463276
rect -6696 459076 590620 459676
rect -4816 455476 588740 456076
rect -2936 451828 586860 452428
rect -8576 444676 592500 445276
rect -6696 441076 590620 441676
rect -4816 437476 588740 438076
rect -2936 433828 586860 434428
rect -8576 426676 592500 427276
rect -6696 423076 590620 423676
rect -4816 419476 588740 420076
rect -2936 415828 586860 416428
rect -8576 408676 592500 409276
rect -6696 405076 590620 405676
rect -4816 401476 588740 402076
rect -2936 397828 586860 398428
rect -8576 390676 592500 391276
rect -6696 387076 590620 387676
rect -4816 383476 588740 384076
rect -2936 379828 586860 380428
rect -8576 372676 592500 373276
rect -6696 369076 590620 369676
rect -4816 365476 588740 366076
rect -2936 361828 586860 362428
rect -8576 354676 592500 355276
rect -6696 351076 590620 351676
rect -4816 347476 588740 348076
rect -2936 343828 586860 344428
rect -8576 336676 592500 337276
rect -6696 333076 590620 333676
rect -4816 329476 588740 330076
rect -2936 325828 586860 326428
rect -8576 318676 592500 319276
rect -6696 315076 590620 315676
rect -4816 311476 588740 312076
rect -2936 307828 586860 308428
rect -8576 300676 592500 301276
rect -6696 297076 590620 297676
rect -4816 293476 588740 294076
rect -2936 289828 586860 290428
rect -8576 282676 592500 283276
rect -6696 279076 590620 279676
rect -4816 275476 588740 276076
rect -2936 271828 586860 272428
rect -8576 264676 592500 265276
rect -6696 261076 590620 261676
rect -4816 257476 588740 258076
rect -2936 253828 586860 254428
rect -8576 246676 592500 247276
rect -6696 243076 590620 243676
rect -4816 239476 588740 240076
rect -2936 235828 586860 236428
rect -8576 228676 592500 229276
rect -6696 225076 590620 225676
rect -4816 221476 588740 222076
rect -2936 217828 586860 218428
rect -8576 210676 592500 211276
rect -6696 207076 590620 207676
rect -4816 203476 588740 204076
rect -2936 199828 586860 200428
rect -8576 192676 592500 193276
rect -6696 189076 590620 189676
rect -4816 185476 588740 186076
rect -2936 181828 586860 182428
rect -8576 174676 592500 175276
rect -6696 171076 590620 171676
rect -4816 167476 588740 168076
rect -2936 163828 586860 164428
rect -8576 156676 592500 157276
rect -6696 153076 590620 153676
rect -4816 149476 588740 150076
rect -2936 145828 586860 146428
rect -8576 138676 592500 139276
rect -6696 135076 590620 135676
rect -4816 131476 588740 132076
rect -2936 127828 586860 128428
rect -8576 120676 592500 121276
rect -6696 117076 590620 117676
rect -4816 113476 588740 114076
rect -2936 109828 586860 110428
rect -8576 102676 592500 103276
rect -6696 99076 590620 99676
rect -4816 95476 588740 96076
rect -2936 91828 586860 92428
rect -8576 84676 592500 85276
rect -6696 81076 590620 81676
rect -4816 77476 588740 78076
rect -2936 73828 586860 74428
rect -8576 66676 592500 67276
rect -6696 63076 590620 63676
rect -4816 59476 588740 60076
rect -2936 55828 586860 56428
rect -8576 48676 592500 49276
rect -6696 45076 590620 45676
rect -4816 41476 588740 42076
rect -2936 37828 586860 38428
rect -8576 30676 592500 31276
rect -6696 27076 590620 27676
rect -4816 23476 588740 24076
rect -2936 19828 586860 20428
rect -8576 12676 592500 13276
rect -6696 9076 590620 9676
rect -4816 5476 588740 6076
rect -2936 1828 586860 2428
rect -1996 -924 585920 -324
rect -2936 -1864 586860 -1264
rect -3876 -2804 587800 -2204
rect -4816 -3744 588740 -3144
rect -5756 -4684 589680 -4084
rect -6696 -5624 590620 -5024
rect -7636 -6564 591560 -5964
rect -8576 -7504 592500 -6904
<< obsm5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect 0 697596 584000 703940
rect -7636 697276 -7036 697278
rect 590960 697276 591560 697278
rect -7636 696674 -7036 696676
rect 590960 696674 591560 696676
rect 0 693996 584000 696356
rect -5756 693676 -5156 693678
rect 589080 693676 589680 693678
rect -5756 693074 -5156 693076
rect 589080 693074 589680 693076
rect 0 690396 584000 692756
rect -3876 690076 -3276 690078
rect 587200 690076 587800 690078
rect -3876 689474 -3276 689476
rect 587200 689474 587800 689476
rect 0 686748 584000 689156
rect -1996 686428 -1396 686430
rect 585320 686428 585920 686430
rect -1996 685826 -1396 685828
rect 585320 685826 585920 685828
rect 0 679596 584000 685508
rect -8576 679276 -7976 679278
rect 591900 679276 592500 679278
rect -8576 678674 -7976 678676
rect 591900 678674 592500 678676
rect 0 675996 584000 678356
rect -6696 675676 -6096 675678
rect 590020 675676 590620 675678
rect -6696 675074 -6096 675076
rect 590020 675074 590620 675076
rect 0 672396 584000 674756
rect -4816 672076 -4216 672078
rect 588140 672076 588740 672078
rect -4816 671474 -4216 671476
rect 588140 671474 588740 671476
rect 0 668748 584000 671156
rect -2936 668428 -2336 668430
rect 586260 668428 586860 668430
rect -2936 667826 -2336 667828
rect 586260 667826 586860 667828
rect 0 661596 584000 667508
rect -7636 661276 -7036 661278
rect 590960 661276 591560 661278
rect -7636 660674 -7036 660676
rect 590960 660674 591560 660676
rect 0 657996 584000 660356
rect -5756 657676 -5156 657678
rect 589080 657676 589680 657678
rect -5756 657074 -5156 657076
rect 589080 657074 589680 657076
rect 0 654396 584000 656756
rect -3876 654076 -3276 654078
rect 587200 654076 587800 654078
rect -3876 653474 -3276 653476
rect 587200 653474 587800 653476
rect 0 650748 584000 653156
rect -1996 650428 -1396 650430
rect 585320 650428 585920 650430
rect -1996 649826 -1396 649828
rect 585320 649826 585920 649828
rect 0 643596 584000 649508
rect -8576 643276 -7976 643278
rect 591900 643276 592500 643278
rect -8576 642674 -7976 642676
rect 591900 642674 592500 642676
rect 0 639996 584000 642356
rect -6696 639676 -6096 639678
rect 590020 639676 590620 639678
rect -6696 639074 -6096 639076
rect 590020 639074 590620 639076
rect 0 636396 584000 638756
rect -4816 636076 -4216 636078
rect 588140 636076 588740 636078
rect -4816 635474 -4216 635476
rect 588140 635474 588740 635476
rect 0 632748 584000 635156
rect -2936 632428 -2336 632430
rect 586260 632428 586860 632430
rect -2936 631826 -2336 631828
rect 586260 631826 586860 631828
rect 0 625596 584000 631508
rect -7636 625276 -7036 625278
rect 590960 625276 591560 625278
rect -7636 624674 -7036 624676
rect 590960 624674 591560 624676
rect 0 621996 584000 624356
rect -5756 621676 -5156 621678
rect 589080 621676 589680 621678
rect -5756 621074 -5156 621076
rect 589080 621074 589680 621076
rect 0 618396 584000 620756
rect -3876 618076 -3276 618078
rect 587200 618076 587800 618078
rect -3876 617474 -3276 617476
rect 587200 617474 587800 617476
rect 0 614748 584000 617156
rect -1996 614428 -1396 614430
rect 585320 614428 585920 614430
rect -1996 613826 -1396 613828
rect 585320 613826 585920 613828
rect 0 607596 584000 613508
rect -8576 607276 -7976 607278
rect 591900 607276 592500 607278
rect -8576 606674 -7976 606676
rect 591900 606674 592500 606676
rect 0 603996 584000 606356
rect -6696 603676 -6096 603678
rect 590020 603676 590620 603678
rect -6696 603074 -6096 603076
rect 590020 603074 590620 603076
rect 0 600396 584000 602756
rect -4816 600076 -4216 600078
rect 588140 600076 588740 600078
rect -4816 599474 -4216 599476
rect 588140 599474 588740 599476
rect 0 596748 584000 599156
rect -2936 596428 -2336 596430
rect 586260 596428 586860 596430
rect -2936 595826 -2336 595828
rect 586260 595826 586860 595828
rect 0 589596 584000 595508
rect -7636 589276 -7036 589278
rect 590960 589276 591560 589278
rect -7636 588674 -7036 588676
rect 590960 588674 591560 588676
rect 0 585996 584000 588356
rect -5756 585676 -5156 585678
rect 589080 585676 589680 585678
rect -5756 585074 -5156 585076
rect 589080 585074 589680 585076
rect 0 582396 584000 584756
rect -3876 582076 -3276 582078
rect 587200 582076 587800 582078
rect -3876 581474 -3276 581476
rect 587200 581474 587800 581476
rect 0 578748 584000 581156
rect -1996 578428 -1396 578430
rect 585320 578428 585920 578430
rect -1996 577826 -1396 577828
rect 585320 577826 585920 577828
rect 0 571596 584000 577508
rect -8576 571276 -7976 571278
rect 591900 571276 592500 571278
rect -8576 570674 -7976 570676
rect 591900 570674 592500 570676
rect 0 567996 584000 570356
rect -6696 567676 -6096 567678
rect 590020 567676 590620 567678
rect -6696 567074 -6096 567076
rect 590020 567074 590620 567076
rect 0 564396 584000 566756
rect -4816 564076 -4216 564078
rect 588140 564076 588740 564078
rect -4816 563474 -4216 563476
rect 588140 563474 588740 563476
rect 0 560748 584000 563156
rect -2936 560428 -2336 560430
rect 586260 560428 586860 560430
rect -2936 559826 -2336 559828
rect 586260 559826 586860 559828
rect 0 553596 584000 559508
rect -7636 553276 -7036 553278
rect 590960 553276 591560 553278
rect -7636 552674 -7036 552676
rect 590960 552674 591560 552676
rect 0 549996 584000 552356
rect -5756 549676 -5156 549678
rect 589080 549676 589680 549678
rect -5756 549074 -5156 549076
rect 589080 549074 589680 549076
rect 0 546396 584000 548756
rect -3876 546076 -3276 546078
rect 587200 546076 587800 546078
rect -3876 545474 -3276 545476
rect 587200 545474 587800 545476
rect 0 542748 584000 545156
rect -1996 542428 -1396 542430
rect 585320 542428 585920 542430
rect -1996 541826 -1396 541828
rect 585320 541826 585920 541828
rect 0 535596 584000 541508
rect -8576 535276 -7976 535278
rect 591900 535276 592500 535278
rect -8576 534674 -7976 534676
rect 591900 534674 592500 534676
rect 0 531996 584000 534356
rect -6696 531676 -6096 531678
rect 590020 531676 590620 531678
rect -6696 531074 -6096 531076
rect 590020 531074 590620 531076
rect 0 528396 584000 530756
rect -4816 528076 -4216 528078
rect 588140 528076 588740 528078
rect -4816 527474 -4216 527476
rect 588140 527474 588740 527476
rect 0 524748 584000 527156
rect -2936 524428 -2336 524430
rect 586260 524428 586860 524430
rect -2936 523826 -2336 523828
rect 586260 523826 586860 523828
rect 0 517596 584000 523508
rect -7636 517276 -7036 517278
rect 590960 517276 591560 517278
rect -7636 516674 -7036 516676
rect 590960 516674 591560 516676
rect 0 513996 584000 516356
rect -5756 513676 -5156 513678
rect 589080 513676 589680 513678
rect -5756 513074 -5156 513076
rect 589080 513074 589680 513076
rect 0 510396 584000 512756
rect -3876 510076 -3276 510078
rect 587200 510076 587800 510078
rect -3876 509474 -3276 509476
rect 587200 509474 587800 509476
rect 0 506748 584000 509156
rect -1996 506428 -1396 506430
rect 585320 506428 585920 506430
rect -1996 505826 -1396 505828
rect 585320 505826 585920 505828
rect 0 499596 584000 505508
rect -8576 499276 -7976 499278
rect 591900 499276 592500 499278
rect -8576 498674 -7976 498676
rect 591900 498674 592500 498676
rect 0 495996 584000 498356
rect -6696 495676 -6096 495678
rect 590020 495676 590620 495678
rect -6696 495074 -6096 495076
rect 590020 495074 590620 495076
rect 0 492396 584000 494756
rect -4816 492076 -4216 492078
rect 588140 492076 588740 492078
rect -4816 491474 -4216 491476
rect 588140 491474 588740 491476
rect 0 488748 584000 491156
rect -2936 488428 -2336 488430
rect 586260 488428 586860 488430
rect -2936 487826 -2336 487828
rect 586260 487826 586860 487828
rect 0 481596 584000 487508
rect -7636 481276 -7036 481278
rect 590960 481276 591560 481278
rect -7636 480674 -7036 480676
rect 590960 480674 591560 480676
rect 0 477996 584000 480356
rect -5756 477676 -5156 477678
rect 589080 477676 589680 477678
rect -5756 477074 -5156 477076
rect 589080 477074 589680 477076
rect 0 474396 584000 476756
rect -3876 474076 -3276 474078
rect 587200 474076 587800 474078
rect -3876 473474 -3276 473476
rect 587200 473474 587800 473476
rect 0 470748 584000 473156
rect -1996 470428 -1396 470430
rect 585320 470428 585920 470430
rect -1996 469826 -1396 469828
rect 585320 469826 585920 469828
rect 0 463596 584000 469508
rect -8576 463276 -7976 463278
rect 591900 463276 592500 463278
rect -8576 462674 -7976 462676
rect 591900 462674 592500 462676
rect 0 459996 584000 462356
rect -6696 459676 -6096 459678
rect 590020 459676 590620 459678
rect -6696 459074 -6096 459076
rect 590020 459074 590620 459076
rect 0 456396 584000 458756
rect -4816 456076 -4216 456078
rect 588140 456076 588740 456078
rect -4816 455474 -4216 455476
rect 588140 455474 588740 455476
rect 0 452748 584000 455156
rect -2936 452428 -2336 452430
rect 586260 452428 586860 452430
rect -2936 451826 -2336 451828
rect 586260 451826 586860 451828
rect 0 445596 584000 451508
rect -7636 445276 -7036 445278
rect 590960 445276 591560 445278
rect -7636 444674 -7036 444676
rect 590960 444674 591560 444676
rect 0 441996 584000 444356
rect -5756 441676 -5156 441678
rect 589080 441676 589680 441678
rect -5756 441074 -5156 441076
rect 589080 441074 589680 441076
rect 0 438396 584000 440756
rect -3876 438076 -3276 438078
rect 587200 438076 587800 438078
rect -3876 437474 -3276 437476
rect 587200 437474 587800 437476
rect 0 434748 584000 437156
rect -1996 434428 -1396 434430
rect 585320 434428 585920 434430
rect -1996 433826 -1396 433828
rect 585320 433826 585920 433828
rect 0 427596 584000 433508
rect -8576 427276 -7976 427278
rect 591900 427276 592500 427278
rect -8576 426674 -7976 426676
rect 591900 426674 592500 426676
rect 0 423996 584000 426356
rect -6696 423676 -6096 423678
rect 590020 423676 590620 423678
rect -6696 423074 -6096 423076
rect 590020 423074 590620 423076
rect 0 420396 584000 422756
rect -4816 420076 -4216 420078
rect 588140 420076 588740 420078
rect -4816 419474 -4216 419476
rect 588140 419474 588740 419476
rect 0 416748 584000 419156
rect -2936 416428 -2336 416430
rect 586260 416428 586860 416430
rect -2936 415826 -2336 415828
rect 586260 415826 586860 415828
rect 0 409596 584000 415508
rect -7636 409276 -7036 409278
rect 590960 409276 591560 409278
rect -7636 408674 -7036 408676
rect 590960 408674 591560 408676
rect 0 405996 584000 408356
rect -5756 405676 -5156 405678
rect 589080 405676 589680 405678
rect -5756 405074 -5156 405076
rect 589080 405074 589680 405076
rect 0 402396 584000 404756
rect -3876 402076 -3276 402078
rect 587200 402076 587800 402078
rect -3876 401474 -3276 401476
rect 587200 401474 587800 401476
rect 0 398748 584000 401156
rect -1996 398428 -1396 398430
rect 585320 398428 585920 398430
rect -1996 397826 -1396 397828
rect 585320 397826 585920 397828
rect 0 391596 584000 397508
rect -8576 391276 -7976 391278
rect 591900 391276 592500 391278
rect -8576 390674 -7976 390676
rect 591900 390674 592500 390676
rect 0 387996 584000 390356
rect -6696 387676 -6096 387678
rect 590020 387676 590620 387678
rect -6696 387074 -6096 387076
rect 590020 387074 590620 387076
rect 0 384396 584000 386756
rect -4816 384076 -4216 384078
rect 588140 384076 588740 384078
rect -4816 383474 -4216 383476
rect 588140 383474 588740 383476
rect 0 380748 584000 383156
rect -2936 380428 -2336 380430
rect 586260 380428 586860 380430
rect -2936 379826 -2336 379828
rect 586260 379826 586860 379828
rect 0 373596 584000 379508
rect -7636 373276 -7036 373278
rect 590960 373276 591560 373278
rect -7636 372674 -7036 372676
rect 590960 372674 591560 372676
rect 0 369996 584000 372356
rect -5756 369676 -5156 369678
rect 589080 369676 589680 369678
rect -5756 369074 -5156 369076
rect 589080 369074 589680 369076
rect 0 366396 584000 368756
rect -3876 366076 -3276 366078
rect 587200 366076 587800 366078
rect -3876 365474 -3276 365476
rect 587200 365474 587800 365476
rect 0 362748 584000 365156
rect -1996 362428 -1396 362430
rect 585320 362428 585920 362430
rect -1996 361826 -1396 361828
rect 585320 361826 585920 361828
rect 0 355596 584000 361508
rect -8576 355276 -7976 355278
rect 591900 355276 592500 355278
rect -8576 354674 -7976 354676
rect 591900 354674 592500 354676
rect 0 351996 584000 354356
rect -6696 351676 -6096 351678
rect 590020 351676 590620 351678
rect -6696 351074 -6096 351076
rect 590020 351074 590620 351076
rect 0 348396 584000 350756
rect -4816 348076 -4216 348078
rect 588140 348076 588740 348078
rect -4816 347474 -4216 347476
rect 588140 347474 588740 347476
rect 0 344748 584000 347156
rect -2936 344428 -2336 344430
rect 586260 344428 586860 344430
rect -2936 343826 -2336 343828
rect 586260 343826 586860 343828
rect 0 337596 584000 343508
rect -7636 337276 -7036 337278
rect 590960 337276 591560 337278
rect -7636 336674 -7036 336676
rect 590960 336674 591560 336676
rect 0 333996 584000 336356
rect -5756 333676 -5156 333678
rect 589080 333676 589680 333678
rect -5756 333074 -5156 333076
rect 589080 333074 589680 333076
rect 0 330396 584000 332756
rect -3876 330076 -3276 330078
rect 587200 330076 587800 330078
rect -3876 329474 -3276 329476
rect 587200 329474 587800 329476
rect 0 326748 584000 329156
rect -1996 326428 -1396 326430
rect 585320 326428 585920 326430
rect -1996 325826 -1396 325828
rect 585320 325826 585920 325828
rect 0 319596 584000 325508
rect -8576 319276 -7976 319278
rect 591900 319276 592500 319278
rect -8576 318674 -7976 318676
rect 591900 318674 592500 318676
rect 0 315996 584000 318356
rect -6696 315676 -6096 315678
rect 590020 315676 590620 315678
rect -6696 315074 -6096 315076
rect 590020 315074 590620 315076
rect 0 312396 584000 314756
rect -4816 312076 -4216 312078
rect 588140 312076 588740 312078
rect -4816 311474 -4216 311476
rect 588140 311474 588740 311476
rect 0 308748 584000 311156
rect -2936 308428 -2336 308430
rect 586260 308428 586860 308430
rect -2936 307826 -2336 307828
rect 586260 307826 586860 307828
rect 0 301596 584000 307508
rect -7636 301276 -7036 301278
rect 590960 301276 591560 301278
rect -7636 300674 -7036 300676
rect 590960 300674 591560 300676
rect 0 297996 584000 300356
rect -5756 297676 -5156 297678
rect 589080 297676 589680 297678
rect -5756 297074 -5156 297076
rect 589080 297074 589680 297076
rect 0 294396 584000 296756
rect -3876 294076 -3276 294078
rect 587200 294076 587800 294078
rect -3876 293474 -3276 293476
rect 587200 293474 587800 293476
rect 0 290748 584000 293156
rect -1996 290428 -1396 290430
rect 585320 290428 585920 290430
rect -1996 289826 -1396 289828
rect 585320 289826 585920 289828
rect 0 283596 584000 289508
rect -8576 283276 -7976 283278
rect 591900 283276 592500 283278
rect -8576 282674 -7976 282676
rect 591900 282674 592500 282676
rect 0 279996 584000 282356
rect -6696 279676 -6096 279678
rect 590020 279676 590620 279678
rect -6696 279074 -6096 279076
rect 590020 279074 590620 279076
rect 0 276396 584000 278756
rect -4816 276076 -4216 276078
rect 588140 276076 588740 276078
rect -4816 275474 -4216 275476
rect 588140 275474 588740 275476
rect 0 272748 584000 275156
rect -2936 272428 -2336 272430
rect 586260 272428 586860 272430
rect -2936 271826 -2336 271828
rect 586260 271826 586860 271828
rect 0 265596 584000 271508
rect -7636 265276 -7036 265278
rect 590960 265276 591560 265278
rect -7636 264674 -7036 264676
rect 590960 264674 591560 264676
rect 0 261996 584000 264356
rect -5756 261676 -5156 261678
rect 589080 261676 589680 261678
rect -5756 261074 -5156 261076
rect 589080 261074 589680 261076
rect 0 258396 584000 260756
rect -3876 258076 -3276 258078
rect 587200 258076 587800 258078
rect -3876 257474 -3276 257476
rect 587200 257474 587800 257476
rect 0 254748 584000 257156
rect -1996 254428 -1396 254430
rect 585320 254428 585920 254430
rect -1996 253826 -1396 253828
rect 585320 253826 585920 253828
rect 0 247596 584000 253508
rect -8576 247276 -7976 247278
rect 591900 247276 592500 247278
rect -8576 246674 -7976 246676
rect 591900 246674 592500 246676
rect 0 243996 584000 246356
rect -6696 243676 -6096 243678
rect 590020 243676 590620 243678
rect -6696 243074 -6096 243076
rect 590020 243074 590620 243076
rect 0 240396 584000 242756
rect -4816 240076 -4216 240078
rect 588140 240076 588740 240078
rect -4816 239474 -4216 239476
rect 588140 239474 588740 239476
rect 0 236748 584000 239156
rect -2936 236428 -2336 236430
rect 586260 236428 586860 236430
rect -2936 235826 -2336 235828
rect 586260 235826 586860 235828
rect 0 229596 584000 235508
rect -7636 229276 -7036 229278
rect 590960 229276 591560 229278
rect -7636 228674 -7036 228676
rect 590960 228674 591560 228676
rect 0 225996 584000 228356
rect -5756 225676 -5156 225678
rect 589080 225676 589680 225678
rect -5756 225074 -5156 225076
rect 589080 225074 589680 225076
rect 0 222396 584000 224756
rect -3876 222076 -3276 222078
rect 587200 222076 587800 222078
rect -3876 221474 -3276 221476
rect 587200 221474 587800 221476
rect 0 218748 584000 221156
rect -1996 218428 -1396 218430
rect 585320 218428 585920 218430
rect -1996 217826 -1396 217828
rect 585320 217826 585920 217828
rect 0 211596 584000 217508
rect -8576 211276 -7976 211278
rect 591900 211276 592500 211278
rect -8576 210674 -7976 210676
rect 591900 210674 592500 210676
rect 0 207996 584000 210356
rect -6696 207676 -6096 207678
rect 590020 207676 590620 207678
rect -6696 207074 -6096 207076
rect 590020 207074 590620 207076
rect 0 204396 584000 206756
rect -4816 204076 -4216 204078
rect 588140 204076 588740 204078
rect -4816 203474 -4216 203476
rect 588140 203474 588740 203476
rect 0 200748 584000 203156
rect -2936 200428 -2336 200430
rect 586260 200428 586860 200430
rect -2936 199826 -2336 199828
rect 586260 199826 586860 199828
rect 0 193596 584000 199508
rect -7636 193276 -7036 193278
rect 590960 193276 591560 193278
rect -7636 192674 -7036 192676
rect 590960 192674 591560 192676
rect 0 189996 584000 192356
rect -5756 189676 -5156 189678
rect 589080 189676 589680 189678
rect -5756 189074 -5156 189076
rect 589080 189074 589680 189076
rect 0 186396 584000 188756
rect -3876 186076 -3276 186078
rect 587200 186076 587800 186078
rect -3876 185474 -3276 185476
rect 587200 185474 587800 185476
rect 0 182748 584000 185156
rect -1996 182428 -1396 182430
rect 585320 182428 585920 182430
rect -1996 181826 -1396 181828
rect 585320 181826 585920 181828
rect 0 175596 584000 181508
rect -8576 175276 -7976 175278
rect 591900 175276 592500 175278
rect -8576 174674 -7976 174676
rect 591900 174674 592500 174676
rect 0 171996 584000 174356
rect -6696 171676 -6096 171678
rect 590020 171676 590620 171678
rect -6696 171074 -6096 171076
rect 590020 171074 590620 171076
rect 0 168396 584000 170756
rect -4816 168076 -4216 168078
rect 588140 168076 588740 168078
rect -4816 167474 -4216 167476
rect 588140 167474 588740 167476
rect 0 164748 584000 167156
rect -2936 164428 -2336 164430
rect 586260 164428 586860 164430
rect -2936 163826 -2336 163828
rect 586260 163826 586860 163828
rect 0 157596 584000 163508
rect -7636 157276 -7036 157278
rect 590960 157276 591560 157278
rect -7636 156674 -7036 156676
rect 590960 156674 591560 156676
rect 0 153996 584000 156356
rect -5756 153676 -5156 153678
rect 589080 153676 589680 153678
rect -5756 153074 -5156 153076
rect 589080 153074 589680 153076
rect 0 150396 584000 152756
rect -3876 150076 -3276 150078
rect 587200 150076 587800 150078
rect -3876 149474 -3276 149476
rect 587200 149474 587800 149476
rect 0 146748 584000 149156
rect -1996 146428 -1396 146430
rect 585320 146428 585920 146430
rect -1996 145826 -1396 145828
rect 585320 145826 585920 145828
rect 0 139596 584000 145508
rect -8576 139276 -7976 139278
rect 591900 139276 592500 139278
rect -8576 138674 -7976 138676
rect 591900 138674 592500 138676
rect 0 135996 584000 138356
rect -6696 135676 -6096 135678
rect 590020 135676 590620 135678
rect -6696 135074 -6096 135076
rect 590020 135074 590620 135076
rect 0 132396 584000 134756
rect -4816 132076 -4216 132078
rect 588140 132076 588740 132078
rect -4816 131474 -4216 131476
rect 588140 131474 588740 131476
rect 0 128748 584000 131156
rect -2936 128428 -2336 128430
rect 586260 128428 586860 128430
rect -2936 127826 -2336 127828
rect 586260 127826 586860 127828
rect 0 121596 584000 127508
rect -7636 121276 -7036 121278
rect 590960 121276 591560 121278
rect -7636 120674 -7036 120676
rect 590960 120674 591560 120676
rect 0 117996 584000 120356
rect -5756 117676 -5156 117678
rect 589080 117676 589680 117678
rect -5756 117074 -5156 117076
rect 589080 117074 589680 117076
rect 0 114396 584000 116756
rect -3876 114076 -3276 114078
rect 587200 114076 587800 114078
rect -3876 113474 -3276 113476
rect 587200 113474 587800 113476
rect 0 110748 584000 113156
rect -1996 110428 -1396 110430
rect 585320 110428 585920 110430
rect -1996 109826 -1396 109828
rect 585320 109826 585920 109828
rect 0 103596 584000 109508
rect -8576 103276 -7976 103278
rect 591900 103276 592500 103278
rect -8576 102674 -7976 102676
rect 591900 102674 592500 102676
rect 0 99996 584000 102356
rect -6696 99676 -6096 99678
rect 590020 99676 590620 99678
rect -6696 99074 -6096 99076
rect 590020 99074 590620 99076
rect 0 96396 584000 98756
rect -4816 96076 -4216 96078
rect 588140 96076 588740 96078
rect -4816 95474 -4216 95476
rect 588140 95474 588740 95476
rect 0 92748 584000 95156
rect -2936 92428 -2336 92430
rect 586260 92428 586860 92430
rect -2936 91826 -2336 91828
rect 586260 91826 586860 91828
rect 0 85596 584000 91508
rect -7636 85276 -7036 85278
rect 590960 85276 591560 85278
rect -7636 84674 -7036 84676
rect 590960 84674 591560 84676
rect 0 81996 584000 84356
rect -5756 81676 -5156 81678
rect 589080 81676 589680 81678
rect -5756 81074 -5156 81076
rect 589080 81074 589680 81076
rect 0 78396 584000 80756
rect -3876 78076 -3276 78078
rect 587200 78076 587800 78078
rect -3876 77474 -3276 77476
rect 587200 77474 587800 77476
rect 0 74748 584000 77156
rect -1996 74428 -1396 74430
rect 585320 74428 585920 74430
rect -1996 73826 -1396 73828
rect 585320 73826 585920 73828
rect 0 67596 584000 73508
rect -8576 67276 -7976 67278
rect 591900 67276 592500 67278
rect -8576 66674 -7976 66676
rect 591900 66674 592500 66676
rect 0 63996 584000 66356
rect -6696 63676 -6096 63678
rect 590020 63676 590620 63678
rect -6696 63074 -6096 63076
rect 590020 63074 590620 63076
rect 0 60396 584000 62756
rect -4816 60076 -4216 60078
rect 588140 60076 588740 60078
rect -4816 59474 -4216 59476
rect 588140 59474 588740 59476
rect 0 56748 584000 59156
rect -2936 56428 -2336 56430
rect 586260 56428 586860 56430
rect -2936 55826 -2336 55828
rect 586260 55826 586860 55828
rect 0 49596 584000 55508
rect -7636 49276 -7036 49278
rect 590960 49276 591560 49278
rect -7636 48674 -7036 48676
rect 590960 48674 591560 48676
rect 0 45996 584000 48356
rect -5756 45676 -5156 45678
rect 589080 45676 589680 45678
rect -5756 45074 -5156 45076
rect 589080 45074 589680 45076
rect 0 42396 584000 44756
rect -3876 42076 -3276 42078
rect 587200 42076 587800 42078
rect -3876 41474 -3276 41476
rect 587200 41474 587800 41476
rect 0 38748 584000 41156
rect -1996 38428 -1396 38430
rect 585320 38428 585920 38430
rect -1996 37826 -1396 37828
rect 585320 37826 585920 37828
rect 0 31596 584000 37508
rect -8576 31276 -7976 31278
rect 591900 31276 592500 31278
rect -8576 30674 -7976 30676
rect 591900 30674 592500 30676
rect 0 27996 584000 30356
rect -6696 27676 -6096 27678
rect 590020 27676 590620 27678
rect -6696 27074 -6096 27076
rect 590020 27074 590620 27076
rect 0 24396 584000 26756
rect -4816 24076 -4216 24078
rect 588140 24076 588740 24078
rect -4816 23474 -4216 23476
rect 588140 23474 588740 23476
rect 0 20748 584000 23156
rect -2936 20428 -2336 20430
rect 586260 20428 586860 20430
rect -2936 19826 -2336 19828
rect 586260 19826 586860 19828
rect 0 13596 584000 19508
rect -7636 13276 -7036 13278
rect 590960 13276 591560 13278
rect -7636 12674 -7036 12676
rect 590960 12674 591560 12676
rect 0 9996 584000 12356
rect -5756 9676 -5156 9678
rect 589080 9676 589680 9678
rect -5756 9074 -5156 9076
rect 589080 9074 589680 9076
rect 0 6396 584000 8756
rect -3876 6076 -3276 6078
rect 587200 6076 587800 6078
rect -3876 5474 -3276 5476
rect 587200 5474 587800 5476
rect 0 2748 584000 5156
rect -1996 2428 -1396 2430
rect 585320 2428 585920 2430
rect -1996 1826 -1396 1828
rect 585320 1826 585920 1828
rect 0 0 584000 1508
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 32 nsew signal input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 33 nsew signal input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 34 nsew signal input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 35 nsew signal input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 36 nsew signal input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 42 nsew signal input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 47 nsew signal input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 48 nsew signal input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 49 nsew signal input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 50 nsew signal input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 51 nsew signal input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 52 nsew signal input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 53 nsew signal input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 54 nsew signal input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 55 nsew signal input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 56 nsew signal input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 57 nsew signal input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 58 nsew signal input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 59 nsew signal input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 60 nsew signal input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 61 nsew signal input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 62 nsew signal input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 63 nsew signal input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 64 nsew signal input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 65 nsew signal input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 66 nsew signal input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 67 nsew signal input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 68 nsew signal input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 69 nsew signal input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 70 nsew signal output
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 71 nsew signal output
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 72 nsew signal output
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 73 nsew signal output
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 74 nsew signal output
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 80 nsew signal output
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 85 nsew signal output
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 86 nsew signal output
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 87 nsew signal output
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 88 nsew signal output
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 89 nsew signal output
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 90 nsew signal output
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 91 nsew signal output
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 92 nsew signal output
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 93 nsew signal output
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 94 nsew signal output
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 95 nsew signal output
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 96 nsew signal output
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 97 nsew signal output
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 98 nsew signal output
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 99 nsew signal output
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 100 nsew signal output
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 101 nsew signal output
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 102 nsew signal output
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 103 nsew signal output
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 104 nsew signal output
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 105 nsew signal output
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 106 nsew signal output
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 107 nsew signal output
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 108 nsew signal output
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 109 nsew signal output
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 110 nsew signal output
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 111 nsew signal output
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 112 nsew signal output
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 118 nsew signal output
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 123 nsew signal output
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 124 nsew signal output
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 125 nsew signal output
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 126 nsew signal output
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 127 nsew signal output
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 128 nsew signal output
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 129 nsew signal output
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 130 nsew signal output
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 131 nsew signal output
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 132 nsew signal output
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 133 nsew signal output
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 134 nsew signal output
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 135 nsew signal output
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 136 nsew signal output
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 137 nsew signal output
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 138 nsew signal output
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 139 nsew signal output
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 140 nsew signal output
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 141 nsew signal output
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 142 nsew signal output
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 143 nsew signal output
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 144 nsew signal output
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 530 nsew signal input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 533 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 599 nsew signal output
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 600 nsew signal output
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 601 nsew signal output
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 602 nsew signal output
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 603 nsew signal output
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 604 nsew signal output
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 605 nsew signal output
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 606 nsew signal output
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 607 nsew signal output
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 608 nsew signal output
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 609 nsew signal output
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 610 nsew signal output
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 611 nsew signal output
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 612 nsew signal output
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 613 nsew signal output
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 614 nsew signal output
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 615 nsew signal output
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 616 nsew signal output
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 617 nsew signal output
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 618 nsew signal output
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 619 nsew signal output
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 620 nsew signal output
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 621 nsew signal output
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 622 nsew signal output
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 623 nsew signal output
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 624 nsew signal output
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 625 nsew signal output
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 626 nsew signal output
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 627 nsew signal output
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 628 nsew signal output
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 629 nsew signal output
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 630 nsew signal output
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 576804 693452 577404 705800 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s 540804 693452 541404 705800 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 504804 693452 505404 705800 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 468804 693452 469404 705800 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 432804 693452 433404 705800 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 396804 693452 397404 705800 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 360804 693452 361404 705800 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 324804 693452 325404 705800 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 288804 693452 289404 705800 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 252804 693452 253404 705800 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 216804 693452 217404 705800 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 180804 693452 181404 705800 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 144804 693452 145404 705800 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 108804 693452 109404 705800 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 72804 693452 73404 705800 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 36804 693452 37404 705800 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 705800 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 654 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 655 nsew power bidirectional
rlabel metal4 s 576804 503452 577404 534548 6 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 540804 503452 541404 534548 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 504804 503452 505404 534548 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 468804 503452 469404 534548 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 432804 503452 433404 534548 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 396804 249452 397404 534548 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 360804 249452 361404 534548 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 324804 -1864 325404 534548 6 vccd1
port 663 nsew power bidirectional
rlabel metal4 s 288804 -1864 289404 534548 6 vccd1
port 664 nsew power bidirectional
rlabel metal4 s 252804 -1864 253404 534548 6 vccd1
port 665 nsew power bidirectional
rlabel metal4 s 216804 249452 217404 534548 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 180804 249452 181404 534548 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 144804 493452 145404 534548 6 vccd1
port 668 nsew power bidirectional
rlabel metal4 s 108804 493452 109404 534548 6 vccd1
port 669 nsew power bidirectional
rlabel metal4 s 72804 493452 73404 534548 6 vccd1
port 670 nsew power bidirectional
rlabel metal4 s 36804 493452 37404 534548 6 vccd1
port 671 nsew power bidirectional
rlabel metal4 s 144804 249452 145404 338548 6 vccd1
port 672 nsew power bidirectional
rlabel metal4 s 108804 249452 109404 338548 6 vccd1
port 673 nsew power bidirectional
rlabel metal4 s 72804 249452 73404 338548 6 vccd1
port 674 nsew power bidirectional
rlabel metal4 s 36804 249452 37404 338548 6 vccd1
port 675 nsew power bidirectional
rlabel metal4 s 576804 249452 577404 334548 6 vccd1
port 676 nsew power bidirectional
rlabel metal4 s 540804 249452 541404 334548 6 vccd1
port 677 nsew power bidirectional
rlabel metal4 s 504804 249452 505404 334548 6 vccd1
port 678 nsew power bidirectional
rlabel metal4 s 468804 249452 469404 334548 6 vccd1
port 679 nsew power bidirectional
rlabel metal4 s 432804 249452 433404 334548 6 vccd1
port 680 nsew power bidirectional
rlabel metal4 s 576804 -1864 577404 10548 6 vccd1
port 681 nsew power bidirectional
rlabel metal4 s 540804 -1864 541404 10548 6 vccd1
port 682 nsew power bidirectional
rlabel metal4 s 504804 -1864 505404 10548 6 vccd1
port 683 nsew power bidirectional
rlabel metal4 s 468804 -1864 469404 10548 6 vccd1
port 684 nsew power bidirectional
rlabel metal4 s 432804 -1864 433404 10548 6 vccd1
port 685 nsew power bidirectional
rlabel metal4 s 396804 -1864 397404 10548 6 vccd1
port 686 nsew power bidirectional
rlabel metal4 s 360804 -1864 361404 10548 6 vccd1
port 687 nsew power bidirectional
rlabel metal4 s 216804 -1864 217404 10548 6 vccd1
port 688 nsew power bidirectional
rlabel metal4 s 180804 -1864 181404 10548 6 vccd1
port 689 nsew power bidirectional
rlabel metal4 s 144804 -1864 145404 10548 6 vccd1
port 690 nsew power bidirectional
rlabel metal4 s 108804 -1864 109404 10548 6 vccd1
port 691 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 10548 6 vccd1
port 692 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 10548 6 vccd1
port 693 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 694 nsew power bidirectional
rlabel metal5 s -2936 685828 586860 686428 6 vccd1
port 695 nsew power bidirectional
rlabel metal5 s -2936 649828 586860 650428 6 vccd1
port 696 nsew power bidirectional
rlabel metal5 s -2936 613828 586860 614428 6 vccd1
port 697 nsew power bidirectional
rlabel metal5 s -2936 577828 586860 578428 6 vccd1
port 698 nsew power bidirectional
rlabel metal5 s -2936 541828 586860 542428 6 vccd1
port 699 nsew power bidirectional
rlabel metal5 s -2936 505828 586860 506428 6 vccd1
port 700 nsew power bidirectional
rlabel metal5 s -2936 469828 586860 470428 6 vccd1
port 701 nsew power bidirectional
rlabel metal5 s -2936 433828 586860 434428 6 vccd1
port 702 nsew power bidirectional
rlabel metal5 s -2936 397828 586860 398428 6 vccd1
port 703 nsew power bidirectional
rlabel metal5 s -2936 361828 586860 362428 6 vccd1
port 704 nsew power bidirectional
rlabel metal5 s -2936 325828 586860 326428 6 vccd1
port 705 nsew power bidirectional
rlabel metal5 s -2936 289828 586860 290428 6 vccd1
port 706 nsew power bidirectional
rlabel metal5 s -2936 253828 586860 254428 6 vccd1
port 707 nsew power bidirectional
rlabel metal5 s -2936 217828 586860 218428 6 vccd1
port 708 nsew power bidirectional
rlabel metal5 s -2936 181828 586860 182428 6 vccd1
port 709 nsew power bidirectional
rlabel metal5 s -2936 145828 586860 146428 6 vccd1
port 710 nsew power bidirectional
rlabel metal5 s -2936 109828 586860 110428 6 vccd1
port 711 nsew power bidirectional
rlabel metal5 s -2936 73828 586860 74428 6 vccd1
port 712 nsew power bidirectional
rlabel metal5 s -2936 37828 586860 38428 6 vccd1
port 713 nsew power bidirectional
rlabel metal5 s -2936 1828 586860 2428 6 vccd1
port 714 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 715 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 716 nsew ground bidirectional
rlabel metal4 s 558804 693452 559404 705800 6 vssd1
port 717 nsew ground bidirectional
rlabel metal4 s 522804 693452 523404 705800 6 vssd1
port 718 nsew ground bidirectional
rlabel metal4 s 486804 693452 487404 705800 6 vssd1
port 719 nsew ground bidirectional
rlabel metal4 s 450804 693452 451404 705800 6 vssd1
port 720 nsew ground bidirectional
rlabel metal4 s 414804 693452 415404 705800 6 vssd1
port 721 nsew ground bidirectional
rlabel metal4 s 378804 693452 379404 705800 6 vssd1
port 722 nsew ground bidirectional
rlabel metal4 s 342804 693452 343404 705800 6 vssd1
port 723 nsew ground bidirectional
rlabel metal4 s 306804 693452 307404 705800 6 vssd1
port 724 nsew ground bidirectional
rlabel metal4 s 270804 693452 271404 705800 6 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 234804 693452 235404 705800 6 vssd1
port 726 nsew ground bidirectional
rlabel metal4 s 198804 693452 199404 705800 6 vssd1
port 727 nsew ground bidirectional
rlabel metal4 s 162804 693452 163404 705800 6 vssd1
port 728 nsew ground bidirectional
rlabel metal4 s 126804 693452 127404 705800 6 vssd1
port 729 nsew ground bidirectional
rlabel metal4 s 90804 693452 91404 705800 6 vssd1
port 730 nsew ground bidirectional
rlabel metal4 s 54804 693452 55404 705800 6 vssd1
port 731 nsew ground bidirectional
rlabel metal4 s 18804 693452 19404 705800 6 vssd1
port 732 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 733 nsew ground bidirectional
rlabel metal4 s 558804 503452 559404 534548 6 vssd1
port 734 nsew ground bidirectional
rlabel metal4 s 522804 503452 523404 534548 6 vssd1
port 735 nsew ground bidirectional
rlabel metal4 s 486804 503452 487404 534548 6 vssd1
port 736 nsew ground bidirectional
rlabel metal4 s 450804 503452 451404 534548 6 vssd1
port 737 nsew ground bidirectional
rlabel metal4 s 414804 503452 415404 534548 6 vssd1
port 738 nsew ground bidirectional
rlabel metal4 s 378804 249452 379404 534548 6 vssd1
port 739 nsew ground bidirectional
rlabel metal4 s 342804 249452 343404 534548 6 vssd1
port 740 nsew ground bidirectional
rlabel metal4 s 306804 -1864 307404 534548 6 vssd1
port 741 nsew ground bidirectional
rlabel metal4 s 270804 -1864 271404 534548 6 vssd1
port 742 nsew ground bidirectional
rlabel metal4 s 234804 249452 235404 534548 6 vssd1
port 743 nsew ground bidirectional
rlabel metal4 s 198804 249452 199404 534548 6 vssd1
port 744 nsew ground bidirectional
rlabel metal4 s 162804 249452 163404 534548 6 vssd1
port 745 nsew ground bidirectional
rlabel metal4 s 126804 493452 127404 534548 6 vssd1
port 746 nsew ground bidirectional
rlabel metal4 s 90804 493452 91404 534548 6 vssd1
port 747 nsew ground bidirectional
rlabel metal4 s 54804 493452 55404 534548 6 vssd1
port 748 nsew ground bidirectional
rlabel metal4 s 18804 493452 19404 534548 6 vssd1
port 749 nsew ground bidirectional
rlabel metal4 s 126804 249452 127404 338548 6 vssd1
port 750 nsew ground bidirectional
rlabel metal4 s 90804 249452 91404 338548 6 vssd1
port 751 nsew ground bidirectional
rlabel metal4 s 54804 249452 55404 338548 6 vssd1
port 752 nsew ground bidirectional
rlabel metal4 s 18804 249452 19404 338548 6 vssd1
port 753 nsew ground bidirectional
rlabel metal4 s 558804 249452 559404 334548 6 vssd1
port 754 nsew ground bidirectional
rlabel metal4 s 522804 249452 523404 334548 6 vssd1
port 755 nsew ground bidirectional
rlabel metal4 s 486804 249452 487404 334548 6 vssd1
port 756 nsew ground bidirectional
rlabel metal4 s 450804 249452 451404 334548 6 vssd1
port 757 nsew ground bidirectional
rlabel metal4 s 414804 249452 415404 334548 6 vssd1
port 758 nsew ground bidirectional
rlabel metal4 s 558804 -1864 559404 10548 6 vssd1
port 759 nsew ground bidirectional
rlabel metal4 s 522804 -1864 523404 10548 6 vssd1
port 760 nsew ground bidirectional
rlabel metal4 s 486804 -1864 487404 10548 6 vssd1
port 761 nsew ground bidirectional
rlabel metal4 s 450804 -1864 451404 10548 6 vssd1
port 762 nsew ground bidirectional
rlabel metal4 s 414804 -1864 415404 10548 6 vssd1
port 763 nsew ground bidirectional
rlabel metal4 s 378804 -1864 379404 10548 6 vssd1
port 764 nsew ground bidirectional
rlabel metal4 s 342804 -1864 343404 10548 6 vssd1
port 765 nsew ground bidirectional
rlabel metal4 s 234804 -1864 235404 10548 6 vssd1
port 766 nsew ground bidirectional
rlabel metal4 s 198804 -1864 199404 10548 6 vssd1
port 767 nsew ground bidirectional
rlabel metal4 s 162804 -1864 163404 10548 6 vssd1
port 768 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 10548 6 vssd1
port 769 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 10548 6 vssd1
port 770 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 10548 6 vssd1
port 771 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 10548 6 vssd1
port 772 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 773 nsew ground bidirectional
rlabel metal5 s -2936 667828 586860 668428 6 vssd1
port 774 nsew ground bidirectional
rlabel metal5 s -2936 631828 586860 632428 6 vssd1
port 775 nsew ground bidirectional
rlabel metal5 s -2936 595828 586860 596428 6 vssd1
port 776 nsew ground bidirectional
rlabel metal5 s -2936 559828 586860 560428 6 vssd1
port 777 nsew ground bidirectional
rlabel metal5 s -2936 523828 586860 524428 6 vssd1
port 778 nsew ground bidirectional
rlabel metal5 s -2936 487828 586860 488428 6 vssd1
port 779 nsew ground bidirectional
rlabel metal5 s -2936 451828 586860 452428 6 vssd1
port 780 nsew ground bidirectional
rlabel metal5 s -2936 415828 586860 416428 6 vssd1
port 781 nsew ground bidirectional
rlabel metal5 s -2936 379828 586860 380428 6 vssd1
port 782 nsew ground bidirectional
rlabel metal5 s -2936 343828 586860 344428 6 vssd1
port 783 nsew ground bidirectional
rlabel metal5 s -2936 307828 586860 308428 6 vssd1
port 784 nsew ground bidirectional
rlabel metal5 s -2936 271828 586860 272428 6 vssd1
port 785 nsew ground bidirectional
rlabel metal5 s -2936 235828 586860 236428 6 vssd1
port 786 nsew ground bidirectional
rlabel metal5 s -2936 199828 586860 200428 6 vssd1
port 787 nsew ground bidirectional
rlabel metal5 s -2936 163828 586860 164428 6 vssd1
port 788 nsew ground bidirectional
rlabel metal5 s -2936 127828 586860 128428 6 vssd1
port 789 nsew ground bidirectional
rlabel metal5 s -2936 91828 586860 92428 6 vssd1
port 790 nsew ground bidirectional
rlabel metal5 s -2936 55828 586860 56428 6 vssd1
port 791 nsew ground bidirectional
rlabel metal5 s -2936 19828 586860 20428 6 vssd1
port 792 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 793 nsew ground bidirectional
rlabel metal4 s 580404 693500 581004 707680 6 vccd2
port 794 nsew power bidirectional
rlabel metal4 s 544404 693500 545004 707680 6 vccd2
port 795 nsew power bidirectional
rlabel metal4 s 508404 693500 509004 707680 6 vccd2
port 796 nsew power bidirectional
rlabel metal4 s 472404 693500 473004 707680 6 vccd2
port 797 nsew power bidirectional
rlabel metal4 s 436404 693500 437004 707680 6 vccd2
port 798 nsew power bidirectional
rlabel metal4 s 400404 693500 401004 707680 6 vccd2
port 799 nsew power bidirectional
rlabel metal4 s 364404 693500 365004 707680 6 vccd2
port 800 nsew power bidirectional
rlabel metal4 s 328404 693500 329004 707680 6 vccd2
port 801 nsew power bidirectional
rlabel metal4 s 292404 693500 293004 707680 6 vccd2
port 802 nsew power bidirectional
rlabel metal4 s 256404 693500 257004 707680 6 vccd2
port 803 nsew power bidirectional
rlabel metal4 s 220404 693500 221004 707680 6 vccd2
port 804 nsew power bidirectional
rlabel metal4 s 184404 693500 185004 707680 6 vccd2
port 805 nsew power bidirectional
rlabel metal4 s 148404 693500 149004 707680 6 vccd2
port 806 nsew power bidirectional
rlabel metal4 s 112404 693500 113004 707680 6 vccd2
port 807 nsew power bidirectional
rlabel metal4 s 76404 693500 77004 707680 6 vccd2
port 808 nsew power bidirectional
rlabel metal4 s 40404 693500 41004 707680 6 vccd2
port 809 nsew power bidirectional
rlabel metal4 s 4404 693500 5004 707680 6 vccd2
port 810 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 811 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 812 nsew power bidirectional
rlabel metal4 s 580404 503500 581004 534500 6 vccd2
port 813 nsew power bidirectional
rlabel metal4 s 544404 503500 545004 534500 6 vccd2
port 814 nsew power bidirectional
rlabel metal4 s 508404 503500 509004 534500 6 vccd2
port 815 nsew power bidirectional
rlabel metal4 s 472404 503500 473004 534500 6 vccd2
port 816 nsew power bidirectional
rlabel metal4 s 436404 503500 437004 534500 6 vccd2
port 817 nsew power bidirectional
rlabel metal4 s 400404 249500 401004 534500 6 vccd2
port 818 nsew power bidirectional
rlabel metal4 s 364404 249500 365004 534500 6 vccd2
port 819 nsew power bidirectional
rlabel metal4 s 328404 -3744 329004 534500 6 vccd2
port 820 nsew power bidirectional
rlabel metal4 s 292404 -3744 293004 534500 6 vccd2
port 821 nsew power bidirectional
rlabel metal4 s 256404 -3744 257004 534500 6 vccd2
port 822 nsew power bidirectional
rlabel metal4 s 220404 249500 221004 534500 6 vccd2
port 823 nsew power bidirectional
rlabel metal4 s 184404 249500 185004 534500 6 vccd2
port 824 nsew power bidirectional
rlabel metal4 s 148404 493500 149004 534500 6 vccd2
port 825 nsew power bidirectional
rlabel metal4 s 112404 493500 113004 534500 6 vccd2
port 826 nsew power bidirectional
rlabel metal4 s 76404 493500 77004 534500 6 vccd2
port 827 nsew power bidirectional
rlabel metal4 s 40404 493500 41004 534500 6 vccd2
port 828 nsew power bidirectional
rlabel metal4 s 4404 493500 5004 534500 6 vccd2
port 829 nsew power bidirectional
rlabel metal4 s 148404 249500 149004 338500 6 vccd2
port 830 nsew power bidirectional
rlabel metal4 s 112404 249500 113004 338500 6 vccd2
port 831 nsew power bidirectional
rlabel metal4 s 76404 249500 77004 338500 6 vccd2
port 832 nsew power bidirectional
rlabel metal4 s 40404 249500 41004 338500 6 vccd2
port 833 nsew power bidirectional
rlabel metal4 s 4404 249500 5004 338500 6 vccd2
port 834 nsew power bidirectional
rlabel metal4 s 580404 249500 581004 334500 6 vccd2
port 835 nsew power bidirectional
rlabel metal4 s 544404 249500 545004 334500 6 vccd2
port 836 nsew power bidirectional
rlabel metal4 s 508404 249500 509004 334500 6 vccd2
port 837 nsew power bidirectional
rlabel metal4 s 472404 249500 473004 334500 6 vccd2
port 838 nsew power bidirectional
rlabel metal4 s 436404 249500 437004 334500 6 vccd2
port 839 nsew power bidirectional
rlabel metal4 s 580404 -3744 581004 10500 6 vccd2
port 840 nsew power bidirectional
rlabel metal4 s 544404 -3744 545004 10500 6 vccd2
port 841 nsew power bidirectional
rlabel metal4 s 508404 -3744 509004 10500 6 vccd2
port 842 nsew power bidirectional
rlabel metal4 s 472404 -3744 473004 10500 6 vccd2
port 843 nsew power bidirectional
rlabel metal4 s 436404 -3744 437004 10500 6 vccd2
port 844 nsew power bidirectional
rlabel metal4 s 400404 -3744 401004 10500 6 vccd2
port 845 nsew power bidirectional
rlabel metal4 s 364404 -3744 365004 10500 6 vccd2
port 846 nsew power bidirectional
rlabel metal4 s 220404 -3744 221004 10500 6 vccd2
port 847 nsew power bidirectional
rlabel metal4 s 184404 -3744 185004 10500 6 vccd2
port 848 nsew power bidirectional
rlabel metal4 s 148404 -3744 149004 10500 6 vccd2
port 849 nsew power bidirectional
rlabel metal4 s 112404 -3744 113004 10500 6 vccd2
port 850 nsew power bidirectional
rlabel metal4 s 76404 -3744 77004 10500 6 vccd2
port 851 nsew power bidirectional
rlabel metal4 s 40404 -3744 41004 10500 6 vccd2
port 852 nsew power bidirectional
rlabel metal4 s 4404 -3744 5004 10500 6 vccd2
port 853 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 854 nsew power bidirectional
rlabel metal5 s -4816 689476 588740 690076 6 vccd2
port 855 nsew power bidirectional
rlabel metal5 s -4816 653476 588740 654076 6 vccd2
port 856 nsew power bidirectional
rlabel metal5 s -4816 617476 588740 618076 6 vccd2
port 857 nsew power bidirectional
rlabel metal5 s -4816 581476 588740 582076 6 vccd2
port 858 nsew power bidirectional
rlabel metal5 s -4816 545476 588740 546076 6 vccd2
port 859 nsew power bidirectional
rlabel metal5 s -4816 509476 588740 510076 6 vccd2
port 860 nsew power bidirectional
rlabel metal5 s -4816 473476 588740 474076 6 vccd2
port 861 nsew power bidirectional
rlabel metal5 s -4816 437476 588740 438076 6 vccd2
port 862 nsew power bidirectional
rlabel metal5 s -4816 401476 588740 402076 6 vccd2
port 863 nsew power bidirectional
rlabel metal5 s -4816 365476 588740 366076 6 vccd2
port 864 nsew power bidirectional
rlabel metal5 s -4816 329476 588740 330076 6 vccd2
port 865 nsew power bidirectional
rlabel metal5 s -4816 293476 588740 294076 6 vccd2
port 866 nsew power bidirectional
rlabel metal5 s -4816 257476 588740 258076 6 vccd2
port 867 nsew power bidirectional
rlabel metal5 s -4816 221476 588740 222076 6 vccd2
port 868 nsew power bidirectional
rlabel metal5 s -4816 185476 588740 186076 6 vccd2
port 869 nsew power bidirectional
rlabel metal5 s -4816 149476 588740 150076 6 vccd2
port 870 nsew power bidirectional
rlabel metal5 s -4816 113476 588740 114076 6 vccd2
port 871 nsew power bidirectional
rlabel metal5 s -4816 77476 588740 78076 6 vccd2
port 872 nsew power bidirectional
rlabel metal5 s -4816 41476 588740 42076 6 vccd2
port 873 nsew power bidirectional
rlabel metal5 s -4816 5476 588740 6076 6 vccd2
port 874 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 875 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 876 nsew ground bidirectional
rlabel metal4 s 562404 693500 563004 707680 6 vssd2
port 877 nsew ground bidirectional
rlabel metal4 s 526404 693500 527004 707680 6 vssd2
port 878 nsew ground bidirectional
rlabel metal4 s 490404 693500 491004 707680 6 vssd2
port 879 nsew ground bidirectional
rlabel metal4 s 454404 693500 455004 707680 6 vssd2
port 880 nsew ground bidirectional
rlabel metal4 s 418404 693500 419004 707680 6 vssd2
port 881 nsew ground bidirectional
rlabel metal4 s 382404 693500 383004 707680 6 vssd2
port 882 nsew ground bidirectional
rlabel metal4 s 346404 693500 347004 707680 6 vssd2
port 883 nsew ground bidirectional
rlabel metal4 s 310404 693500 311004 707680 6 vssd2
port 884 nsew ground bidirectional
rlabel metal4 s 274404 693500 275004 707680 6 vssd2
port 885 nsew ground bidirectional
rlabel metal4 s 238404 693500 239004 707680 6 vssd2
port 886 nsew ground bidirectional
rlabel metal4 s 202404 693500 203004 707680 6 vssd2
port 887 nsew ground bidirectional
rlabel metal4 s 166404 693500 167004 707680 6 vssd2
port 888 nsew ground bidirectional
rlabel metal4 s 130404 693500 131004 707680 6 vssd2
port 889 nsew ground bidirectional
rlabel metal4 s 94404 693500 95004 707680 6 vssd2
port 890 nsew ground bidirectional
rlabel metal4 s 58404 693500 59004 707680 6 vssd2
port 891 nsew ground bidirectional
rlabel metal4 s 22404 693500 23004 707680 6 vssd2
port 892 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 893 nsew ground bidirectional
rlabel metal4 s 562404 503500 563004 534500 6 vssd2
port 894 nsew ground bidirectional
rlabel metal4 s 526404 503500 527004 534500 6 vssd2
port 895 nsew ground bidirectional
rlabel metal4 s 490404 503500 491004 534500 6 vssd2
port 896 nsew ground bidirectional
rlabel metal4 s 454404 503500 455004 534500 6 vssd2
port 897 nsew ground bidirectional
rlabel metal4 s 418404 503500 419004 534500 6 vssd2
port 898 nsew ground bidirectional
rlabel metal4 s 382404 249500 383004 534500 6 vssd2
port 899 nsew ground bidirectional
rlabel metal4 s 346404 249500 347004 534500 6 vssd2
port 900 nsew ground bidirectional
rlabel metal4 s 310404 -3744 311004 534500 6 vssd2
port 901 nsew ground bidirectional
rlabel metal4 s 274404 -3744 275004 534500 6 vssd2
port 902 nsew ground bidirectional
rlabel metal4 s 238404 249500 239004 534500 6 vssd2
port 903 nsew ground bidirectional
rlabel metal4 s 202404 249500 203004 534500 6 vssd2
port 904 nsew ground bidirectional
rlabel metal4 s 166404 249500 167004 534500 6 vssd2
port 905 nsew ground bidirectional
rlabel metal4 s 130404 493500 131004 534500 6 vssd2
port 906 nsew ground bidirectional
rlabel metal4 s 94404 493500 95004 534500 6 vssd2
port 907 nsew ground bidirectional
rlabel metal4 s 58404 493500 59004 534500 6 vssd2
port 908 nsew ground bidirectional
rlabel metal4 s 22404 493500 23004 534500 6 vssd2
port 909 nsew ground bidirectional
rlabel metal4 s 130404 249500 131004 338500 6 vssd2
port 910 nsew ground bidirectional
rlabel metal4 s 94404 249500 95004 338500 6 vssd2
port 911 nsew ground bidirectional
rlabel metal4 s 58404 249500 59004 338500 6 vssd2
port 912 nsew ground bidirectional
rlabel metal4 s 22404 249500 23004 338500 6 vssd2
port 913 nsew ground bidirectional
rlabel metal4 s 562404 249500 563004 334500 6 vssd2
port 914 nsew ground bidirectional
rlabel metal4 s 526404 249500 527004 334500 6 vssd2
port 915 nsew ground bidirectional
rlabel metal4 s 490404 249500 491004 334500 6 vssd2
port 916 nsew ground bidirectional
rlabel metal4 s 454404 249500 455004 334500 6 vssd2
port 917 nsew ground bidirectional
rlabel metal4 s 418404 249500 419004 334500 6 vssd2
port 918 nsew ground bidirectional
rlabel metal4 s 562404 -3744 563004 10500 6 vssd2
port 919 nsew ground bidirectional
rlabel metal4 s 526404 -3744 527004 10500 6 vssd2
port 920 nsew ground bidirectional
rlabel metal4 s 490404 -3744 491004 10500 6 vssd2
port 921 nsew ground bidirectional
rlabel metal4 s 454404 -3744 455004 10500 6 vssd2
port 922 nsew ground bidirectional
rlabel metal4 s 418404 -3744 419004 10500 6 vssd2
port 923 nsew ground bidirectional
rlabel metal4 s 382404 -3744 383004 10500 6 vssd2
port 924 nsew ground bidirectional
rlabel metal4 s 346404 -3744 347004 10500 6 vssd2
port 925 nsew ground bidirectional
rlabel metal4 s 238404 -3744 239004 10500 6 vssd2
port 926 nsew ground bidirectional
rlabel metal4 s 202404 -3744 203004 10500 6 vssd2
port 927 nsew ground bidirectional
rlabel metal4 s 166404 -3744 167004 10500 6 vssd2
port 928 nsew ground bidirectional
rlabel metal4 s 130404 -3744 131004 10500 6 vssd2
port 929 nsew ground bidirectional
rlabel metal4 s 94404 -3744 95004 10500 6 vssd2
port 930 nsew ground bidirectional
rlabel metal4 s 58404 -3744 59004 10500 6 vssd2
port 931 nsew ground bidirectional
rlabel metal4 s 22404 -3744 23004 10500 6 vssd2
port 932 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 933 nsew ground bidirectional
rlabel metal5 s -4816 671476 588740 672076 6 vssd2
port 934 nsew ground bidirectional
rlabel metal5 s -4816 635476 588740 636076 6 vssd2
port 935 nsew ground bidirectional
rlabel metal5 s -4816 599476 588740 600076 6 vssd2
port 936 nsew ground bidirectional
rlabel metal5 s -4816 563476 588740 564076 6 vssd2
port 937 nsew ground bidirectional
rlabel metal5 s -4816 527476 588740 528076 6 vssd2
port 938 nsew ground bidirectional
rlabel metal5 s -4816 491476 588740 492076 6 vssd2
port 939 nsew ground bidirectional
rlabel metal5 s -4816 455476 588740 456076 6 vssd2
port 940 nsew ground bidirectional
rlabel metal5 s -4816 419476 588740 420076 6 vssd2
port 941 nsew ground bidirectional
rlabel metal5 s -4816 383476 588740 384076 6 vssd2
port 942 nsew ground bidirectional
rlabel metal5 s -4816 347476 588740 348076 6 vssd2
port 943 nsew ground bidirectional
rlabel metal5 s -4816 311476 588740 312076 6 vssd2
port 944 nsew ground bidirectional
rlabel metal5 s -4816 275476 588740 276076 6 vssd2
port 945 nsew ground bidirectional
rlabel metal5 s -4816 239476 588740 240076 6 vssd2
port 946 nsew ground bidirectional
rlabel metal5 s -4816 203476 588740 204076 6 vssd2
port 947 nsew ground bidirectional
rlabel metal5 s -4816 167476 588740 168076 6 vssd2
port 948 nsew ground bidirectional
rlabel metal5 s -4816 131476 588740 132076 6 vssd2
port 949 nsew ground bidirectional
rlabel metal5 s -4816 95476 588740 96076 6 vssd2
port 950 nsew ground bidirectional
rlabel metal5 s -4816 59476 588740 60076 6 vssd2
port 951 nsew ground bidirectional
rlabel metal5 s -4816 23476 588740 24076 6 vssd2
port 952 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 953 nsew ground bidirectional
rlabel metal4 s 548004 693500 548604 709560 6 vdda1
port 954 nsew power bidirectional
rlabel metal4 s 512004 693500 512604 709560 6 vdda1
port 955 nsew power bidirectional
rlabel metal4 s 476004 693500 476604 709560 6 vdda1
port 956 nsew power bidirectional
rlabel metal4 s 440004 693500 440604 709560 6 vdda1
port 957 nsew power bidirectional
rlabel metal4 s 404004 693500 404604 709560 6 vdda1
port 958 nsew power bidirectional
rlabel metal4 s 368004 693500 368604 709560 6 vdda1
port 959 nsew power bidirectional
rlabel metal4 s 332004 693500 332604 709560 6 vdda1
port 960 nsew power bidirectional
rlabel metal4 s 296004 693500 296604 709560 6 vdda1
port 961 nsew power bidirectional
rlabel metal4 s 260004 693500 260604 709560 6 vdda1
port 962 nsew power bidirectional
rlabel metal4 s 224004 693500 224604 709560 6 vdda1
port 963 nsew power bidirectional
rlabel metal4 s 188004 693500 188604 709560 6 vdda1
port 964 nsew power bidirectional
rlabel metal4 s 152004 693500 152604 709560 6 vdda1
port 965 nsew power bidirectional
rlabel metal4 s 116004 693500 116604 709560 6 vdda1
port 966 nsew power bidirectional
rlabel metal4 s 80004 693500 80604 709560 6 vdda1
port 967 nsew power bidirectional
rlabel metal4 s 44004 693500 44604 709560 6 vdda1
port 968 nsew power bidirectional
rlabel metal4 s 8004 693500 8604 709560 6 vdda1
port 969 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 970 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 971 nsew power bidirectional
rlabel metal4 s 548004 503500 548604 534500 6 vdda1
port 972 nsew power bidirectional
rlabel metal4 s 512004 503500 512604 534500 6 vdda1
port 973 nsew power bidirectional
rlabel metal4 s 476004 503500 476604 534500 6 vdda1
port 974 nsew power bidirectional
rlabel metal4 s 440004 503500 440604 534500 6 vdda1
port 975 nsew power bidirectional
rlabel metal4 s 404004 249500 404604 534500 6 vdda1
port 976 nsew power bidirectional
rlabel metal4 s 368004 249500 368604 534500 6 vdda1
port 977 nsew power bidirectional
rlabel metal4 s 332004 -5624 332604 534500 6 vdda1
port 978 nsew power bidirectional
rlabel metal4 s 296004 -5624 296604 534500 6 vdda1
port 979 nsew power bidirectional
rlabel metal4 s 260004 -5624 260604 534500 6 vdda1
port 980 nsew power bidirectional
rlabel metal4 s 224004 249500 224604 534500 6 vdda1
port 981 nsew power bidirectional
rlabel metal4 s 188004 249500 188604 534500 6 vdda1
port 982 nsew power bidirectional
rlabel metal4 s 152004 493500 152604 534500 6 vdda1
port 983 nsew power bidirectional
rlabel metal4 s 116004 493500 116604 534500 6 vdda1
port 984 nsew power bidirectional
rlabel metal4 s 80004 493500 80604 534500 6 vdda1
port 985 nsew power bidirectional
rlabel metal4 s 44004 493500 44604 534500 6 vdda1
port 986 nsew power bidirectional
rlabel metal4 s 8004 493500 8604 534500 6 vdda1
port 987 nsew power bidirectional
rlabel metal4 s 152004 249500 152604 338500 6 vdda1
port 988 nsew power bidirectional
rlabel metal4 s 116004 249500 116604 338500 6 vdda1
port 989 nsew power bidirectional
rlabel metal4 s 80004 249500 80604 338500 6 vdda1
port 990 nsew power bidirectional
rlabel metal4 s 44004 249500 44604 338500 6 vdda1
port 991 nsew power bidirectional
rlabel metal4 s 8004 249500 8604 338500 6 vdda1
port 992 nsew power bidirectional
rlabel metal4 s 548004 249500 548604 334500 6 vdda1
port 993 nsew power bidirectional
rlabel metal4 s 512004 249500 512604 334500 6 vdda1
port 994 nsew power bidirectional
rlabel metal4 s 476004 249500 476604 334500 6 vdda1
port 995 nsew power bidirectional
rlabel metal4 s 440004 249500 440604 334500 6 vdda1
port 996 nsew power bidirectional
rlabel metal4 s 548004 -5624 548604 10500 6 vdda1
port 997 nsew power bidirectional
rlabel metal4 s 512004 -5624 512604 10500 6 vdda1
port 998 nsew power bidirectional
rlabel metal4 s 476004 -5624 476604 10500 6 vdda1
port 999 nsew power bidirectional
rlabel metal4 s 440004 -5624 440604 10500 6 vdda1
port 1000 nsew power bidirectional
rlabel metal4 s 404004 -5624 404604 10500 6 vdda1
port 1001 nsew power bidirectional
rlabel metal4 s 368004 -5624 368604 10500 6 vdda1
port 1002 nsew power bidirectional
rlabel metal4 s 224004 -5624 224604 10500 6 vdda1
port 1003 nsew power bidirectional
rlabel metal4 s 188004 -5624 188604 10500 6 vdda1
port 1004 nsew power bidirectional
rlabel metal4 s 152004 -5624 152604 10500 6 vdda1
port 1005 nsew power bidirectional
rlabel metal4 s 116004 -5624 116604 10500 6 vdda1
port 1006 nsew power bidirectional
rlabel metal4 s 80004 -5624 80604 10500 6 vdda1
port 1007 nsew power bidirectional
rlabel metal4 s 44004 -5624 44604 10500 6 vdda1
port 1008 nsew power bidirectional
rlabel metal4 s 8004 -5624 8604 10500 6 vdda1
port 1009 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 1010 nsew power bidirectional
rlabel metal5 s -6696 693076 590620 693676 6 vdda1
port 1011 nsew power bidirectional
rlabel metal5 s -6696 657076 590620 657676 6 vdda1
port 1012 nsew power bidirectional
rlabel metal5 s -6696 621076 590620 621676 6 vdda1
port 1013 nsew power bidirectional
rlabel metal5 s -6696 585076 590620 585676 6 vdda1
port 1014 nsew power bidirectional
rlabel metal5 s -6696 549076 590620 549676 6 vdda1
port 1015 nsew power bidirectional
rlabel metal5 s -6696 513076 590620 513676 6 vdda1
port 1016 nsew power bidirectional
rlabel metal5 s -6696 477076 590620 477676 6 vdda1
port 1017 nsew power bidirectional
rlabel metal5 s -6696 441076 590620 441676 6 vdda1
port 1018 nsew power bidirectional
rlabel metal5 s -6696 405076 590620 405676 6 vdda1
port 1019 nsew power bidirectional
rlabel metal5 s -6696 369076 590620 369676 6 vdda1
port 1020 nsew power bidirectional
rlabel metal5 s -6696 333076 590620 333676 6 vdda1
port 1021 nsew power bidirectional
rlabel metal5 s -6696 297076 590620 297676 6 vdda1
port 1022 nsew power bidirectional
rlabel metal5 s -6696 261076 590620 261676 6 vdda1
port 1023 nsew power bidirectional
rlabel metal5 s -6696 225076 590620 225676 6 vdda1
port 1024 nsew power bidirectional
rlabel metal5 s -6696 189076 590620 189676 6 vdda1
port 1025 nsew power bidirectional
rlabel metal5 s -6696 153076 590620 153676 6 vdda1
port 1026 nsew power bidirectional
rlabel metal5 s -6696 117076 590620 117676 6 vdda1
port 1027 nsew power bidirectional
rlabel metal5 s -6696 81076 590620 81676 6 vdda1
port 1028 nsew power bidirectional
rlabel metal5 s -6696 45076 590620 45676 6 vdda1
port 1029 nsew power bidirectional
rlabel metal5 s -6696 9076 590620 9676 6 vdda1
port 1030 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 1031 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 1032 nsew ground bidirectional
rlabel metal4 s 566004 693500 566604 709560 6 vssa1
port 1033 nsew ground bidirectional
rlabel metal4 s 530004 693500 530604 709560 6 vssa1
port 1034 nsew ground bidirectional
rlabel metal4 s 494004 693500 494604 709560 6 vssa1
port 1035 nsew ground bidirectional
rlabel metal4 s 458004 693500 458604 709560 6 vssa1
port 1036 nsew ground bidirectional
rlabel metal4 s 422004 693500 422604 709560 6 vssa1
port 1037 nsew ground bidirectional
rlabel metal4 s 386004 693500 386604 709560 6 vssa1
port 1038 nsew ground bidirectional
rlabel metal4 s 350004 693500 350604 709560 6 vssa1
port 1039 nsew ground bidirectional
rlabel metal4 s 314004 693500 314604 709560 6 vssa1
port 1040 nsew ground bidirectional
rlabel metal4 s 278004 693500 278604 709560 6 vssa1
port 1041 nsew ground bidirectional
rlabel metal4 s 242004 693500 242604 709560 6 vssa1
port 1042 nsew ground bidirectional
rlabel metal4 s 206004 693500 206604 709560 6 vssa1
port 1043 nsew ground bidirectional
rlabel metal4 s 170004 693500 170604 709560 6 vssa1
port 1044 nsew ground bidirectional
rlabel metal4 s 134004 693500 134604 709560 6 vssa1
port 1045 nsew ground bidirectional
rlabel metal4 s 98004 693500 98604 709560 6 vssa1
port 1046 nsew ground bidirectional
rlabel metal4 s 62004 693500 62604 709560 6 vssa1
port 1047 nsew ground bidirectional
rlabel metal4 s 26004 693500 26604 709560 6 vssa1
port 1048 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 1049 nsew ground bidirectional
rlabel metal4 s 566004 503500 566604 534500 6 vssa1
port 1050 nsew ground bidirectional
rlabel metal4 s 530004 503500 530604 534500 6 vssa1
port 1051 nsew ground bidirectional
rlabel metal4 s 494004 503500 494604 534500 6 vssa1
port 1052 nsew ground bidirectional
rlabel metal4 s 458004 503500 458604 534500 6 vssa1
port 1053 nsew ground bidirectional
rlabel metal4 s 422004 503500 422604 534500 6 vssa1
port 1054 nsew ground bidirectional
rlabel metal4 s 386004 249500 386604 534500 6 vssa1
port 1055 nsew ground bidirectional
rlabel metal4 s 350004 249500 350604 534500 6 vssa1
port 1056 nsew ground bidirectional
rlabel metal4 s 314004 -5624 314604 534500 6 vssa1
port 1057 nsew ground bidirectional
rlabel metal4 s 278004 -5624 278604 534500 6 vssa1
port 1058 nsew ground bidirectional
rlabel metal4 s 242004 -5624 242604 534500 6 vssa1
port 1059 nsew ground bidirectional
rlabel metal4 s 206004 249500 206604 534500 6 vssa1
port 1060 nsew ground bidirectional
rlabel metal4 s 170004 249500 170604 534500 6 vssa1
port 1061 nsew ground bidirectional
rlabel metal4 s 134004 493500 134604 534500 6 vssa1
port 1062 nsew ground bidirectional
rlabel metal4 s 98004 493500 98604 534500 6 vssa1
port 1063 nsew ground bidirectional
rlabel metal4 s 62004 493500 62604 534500 6 vssa1
port 1064 nsew ground bidirectional
rlabel metal4 s 26004 493500 26604 534500 6 vssa1
port 1065 nsew ground bidirectional
rlabel metal4 s 134004 249500 134604 338500 6 vssa1
port 1066 nsew ground bidirectional
rlabel metal4 s 98004 249500 98604 338500 6 vssa1
port 1067 nsew ground bidirectional
rlabel metal4 s 62004 249500 62604 338500 6 vssa1
port 1068 nsew ground bidirectional
rlabel metal4 s 26004 249500 26604 338500 6 vssa1
port 1069 nsew ground bidirectional
rlabel metal4 s 566004 249500 566604 334500 6 vssa1
port 1070 nsew ground bidirectional
rlabel metal4 s 530004 249500 530604 334500 6 vssa1
port 1071 nsew ground bidirectional
rlabel metal4 s 494004 249500 494604 334500 6 vssa1
port 1072 nsew ground bidirectional
rlabel metal4 s 458004 249500 458604 334500 6 vssa1
port 1073 nsew ground bidirectional
rlabel metal4 s 422004 249500 422604 334500 6 vssa1
port 1074 nsew ground bidirectional
rlabel metal4 s 566004 -5624 566604 10500 6 vssa1
port 1075 nsew ground bidirectional
rlabel metal4 s 530004 -5624 530604 10500 6 vssa1
port 1076 nsew ground bidirectional
rlabel metal4 s 494004 -5624 494604 10500 6 vssa1
port 1077 nsew ground bidirectional
rlabel metal4 s 458004 -5624 458604 10500 6 vssa1
port 1078 nsew ground bidirectional
rlabel metal4 s 422004 -5624 422604 10500 6 vssa1
port 1079 nsew ground bidirectional
rlabel metal4 s 386004 -5624 386604 10500 6 vssa1
port 1080 nsew ground bidirectional
rlabel metal4 s 350004 -5624 350604 10500 6 vssa1
port 1081 nsew ground bidirectional
rlabel metal4 s 206004 -5624 206604 10500 6 vssa1
port 1082 nsew ground bidirectional
rlabel metal4 s 170004 -5624 170604 10500 6 vssa1
port 1083 nsew ground bidirectional
rlabel metal4 s 134004 -5624 134604 10500 6 vssa1
port 1084 nsew ground bidirectional
rlabel metal4 s 98004 -5624 98604 10500 6 vssa1
port 1085 nsew ground bidirectional
rlabel metal4 s 62004 -5624 62604 10500 6 vssa1
port 1086 nsew ground bidirectional
rlabel metal4 s 26004 -5624 26604 10500 6 vssa1
port 1087 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 1088 nsew ground bidirectional
rlabel metal5 s -6696 675076 590620 675676 6 vssa1
port 1089 nsew ground bidirectional
rlabel metal5 s -6696 639076 590620 639676 6 vssa1
port 1090 nsew ground bidirectional
rlabel metal5 s -6696 603076 590620 603676 6 vssa1
port 1091 nsew ground bidirectional
rlabel metal5 s -6696 567076 590620 567676 6 vssa1
port 1092 nsew ground bidirectional
rlabel metal5 s -6696 531076 590620 531676 6 vssa1
port 1093 nsew ground bidirectional
rlabel metal5 s -6696 495076 590620 495676 6 vssa1
port 1094 nsew ground bidirectional
rlabel metal5 s -6696 459076 590620 459676 6 vssa1
port 1095 nsew ground bidirectional
rlabel metal5 s -6696 423076 590620 423676 6 vssa1
port 1096 nsew ground bidirectional
rlabel metal5 s -6696 387076 590620 387676 6 vssa1
port 1097 nsew ground bidirectional
rlabel metal5 s -6696 351076 590620 351676 6 vssa1
port 1098 nsew ground bidirectional
rlabel metal5 s -6696 315076 590620 315676 6 vssa1
port 1099 nsew ground bidirectional
rlabel metal5 s -6696 279076 590620 279676 6 vssa1
port 1100 nsew ground bidirectional
rlabel metal5 s -6696 243076 590620 243676 6 vssa1
port 1101 nsew ground bidirectional
rlabel metal5 s -6696 207076 590620 207676 6 vssa1
port 1102 nsew ground bidirectional
rlabel metal5 s -6696 171076 590620 171676 6 vssa1
port 1103 nsew ground bidirectional
rlabel metal5 s -6696 135076 590620 135676 6 vssa1
port 1104 nsew ground bidirectional
rlabel metal5 s -6696 99076 590620 99676 6 vssa1
port 1105 nsew ground bidirectional
rlabel metal5 s -6696 63076 590620 63676 6 vssa1
port 1106 nsew ground bidirectional
rlabel metal5 s -6696 27076 590620 27676 6 vssa1
port 1107 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 1108 nsew ground bidirectional
rlabel metal4 s 551604 693500 552204 711440 6 vdda2
port 1109 nsew power bidirectional
rlabel metal4 s 515604 693500 516204 711440 6 vdda2
port 1110 nsew power bidirectional
rlabel metal4 s 479604 693500 480204 711440 6 vdda2
port 1111 nsew power bidirectional
rlabel metal4 s 443604 693500 444204 711440 6 vdda2
port 1112 nsew power bidirectional
rlabel metal4 s 407604 693500 408204 711440 6 vdda2
port 1113 nsew power bidirectional
rlabel metal4 s 371604 693500 372204 711440 6 vdda2
port 1114 nsew power bidirectional
rlabel metal4 s 335604 693500 336204 711440 6 vdda2
port 1115 nsew power bidirectional
rlabel metal4 s 299604 693500 300204 711440 6 vdda2
port 1116 nsew power bidirectional
rlabel metal4 s 263604 693500 264204 711440 6 vdda2
port 1117 nsew power bidirectional
rlabel metal4 s 227604 693500 228204 711440 6 vdda2
port 1118 nsew power bidirectional
rlabel metal4 s 191604 693500 192204 711440 6 vdda2
port 1119 nsew power bidirectional
rlabel metal4 s 155604 693500 156204 711440 6 vdda2
port 1120 nsew power bidirectional
rlabel metal4 s 119604 693500 120204 711440 6 vdda2
port 1121 nsew power bidirectional
rlabel metal4 s 83604 693500 84204 711440 6 vdda2
port 1122 nsew power bidirectional
rlabel metal4 s 47604 693500 48204 711440 6 vdda2
port 1123 nsew power bidirectional
rlabel metal4 s 11604 693500 12204 711440 6 vdda2
port 1124 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 1125 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 1126 nsew power bidirectional
rlabel metal4 s 551604 503500 552204 534500 6 vdda2
port 1127 nsew power bidirectional
rlabel metal4 s 515604 503500 516204 534500 6 vdda2
port 1128 nsew power bidirectional
rlabel metal4 s 479604 503500 480204 534500 6 vdda2
port 1129 nsew power bidirectional
rlabel metal4 s 443604 503500 444204 534500 6 vdda2
port 1130 nsew power bidirectional
rlabel metal4 s 407604 249500 408204 534500 6 vdda2
port 1131 nsew power bidirectional
rlabel metal4 s 371604 249500 372204 534500 6 vdda2
port 1132 nsew power bidirectional
rlabel metal4 s 335604 -7504 336204 534500 6 vdda2
port 1133 nsew power bidirectional
rlabel metal4 s 299604 -7504 300204 534500 6 vdda2
port 1134 nsew power bidirectional
rlabel metal4 s 263604 -7504 264204 534500 6 vdda2
port 1135 nsew power bidirectional
rlabel metal4 s 227604 249500 228204 534500 6 vdda2
port 1136 nsew power bidirectional
rlabel metal4 s 191604 249500 192204 534500 6 vdda2
port 1137 nsew power bidirectional
rlabel metal4 s 155604 493500 156204 534500 6 vdda2
port 1138 nsew power bidirectional
rlabel metal4 s 119604 493500 120204 534500 6 vdda2
port 1139 nsew power bidirectional
rlabel metal4 s 83604 493500 84204 534500 6 vdda2
port 1140 nsew power bidirectional
rlabel metal4 s 47604 493500 48204 534500 6 vdda2
port 1141 nsew power bidirectional
rlabel metal4 s 11604 493500 12204 534500 6 vdda2
port 1142 nsew power bidirectional
rlabel metal4 s 155604 249500 156204 338500 6 vdda2
port 1143 nsew power bidirectional
rlabel metal4 s 119604 249500 120204 338500 6 vdda2
port 1144 nsew power bidirectional
rlabel metal4 s 83604 249500 84204 338500 6 vdda2
port 1145 nsew power bidirectional
rlabel metal4 s 47604 249500 48204 338500 6 vdda2
port 1146 nsew power bidirectional
rlabel metal4 s 11604 249500 12204 338500 6 vdda2
port 1147 nsew power bidirectional
rlabel metal4 s 551604 249500 552204 334500 6 vdda2
port 1148 nsew power bidirectional
rlabel metal4 s 515604 249500 516204 334500 6 vdda2
port 1149 nsew power bidirectional
rlabel metal4 s 479604 249500 480204 334500 6 vdda2
port 1150 nsew power bidirectional
rlabel metal4 s 443604 249500 444204 334500 6 vdda2
port 1151 nsew power bidirectional
rlabel metal4 s 551604 -7504 552204 10500 6 vdda2
port 1152 nsew power bidirectional
rlabel metal4 s 515604 -7504 516204 10500 6 vdda2
port 1153 nsew power bidirectional
rlabel metal4 s 479604 -7504 480204 10500 6 vdda2
port 1154 nsew power bidirectional
rlabel metal4 s 443604 -7504 444204 10500 6 vdda2
port 1155 nsew power bidirectional
rlabel metal4 s 407604 -7504 408204 10500 6 vdda2
port 1156 nsew power bidirectional
rlabel metal4 s 371604 -7504 372204 10500 6 vdda2
port 1157 nsew power bidirectional
rlabel metal4 s 227604 -7504 228204 10500 6 vdda2
port 1158 nsew power bidirectional
rlabel metal4 s 191604 -7504 192204 10500 6 vdda2
port 1159 nsew power bidirectional
rlabel metal4 s 155604 -7504 156204 10500 6 vdda2
port 1160 nsew power bidirectional
rlabel metal4 s 119604 -7504 120204 10500 6 vdda2
port 1161 nsew power bidirectional
rlabel metal4 s 83604 -7504 84204 10500 6 vdda2
port 1162 nsew power bidirectional
rlabel metal4 s 47604 -7504 48204 10500 6 vdda2
port 1163 nsew power bidirectional
rlabel metal4 s 11604 -7504 12204 10500 6 vdda2
port 1164 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 1165 nsew power bidirectional
rlabel metal5 s -8576 696676 592500 697276 6 vdda2
port 1166 nsew power bidirectional
rlabel metal5 s -8576 660676 592500 661276 6 vdda2
port 1167 nsew power bidirectional
rlabel metal5 s -8576 624676 592500 625276 6 vdda2
port 1168 nsew power bidirectional
rlabel metal5 s -8576 588676 592500 589276 6 vdda2
port 1169 nsew power bidirectional
rlabel metal5 s -8576 552676 592500 553276 6 vdda2
port 1170 nsew power bidirectional
rlabel metal5 s -8576 516676 592500 517276 6 vdda2
port 1171 nsew power bidirectional
rlabel metal5 s -8576 480676 592500 481276 6 vdda2
port 1172 nsew power bidirectional
rlabel metal5 s -8576 444676 592500 445276 6 vdda2
port 1173 nsew power bidirectional
rlabel metal5 s -8576 408676 592500 409276 6 vdda2
port 1174 nsew power bidirectional
rlabel metal5 s -8576 372676 592500 373276 6 vdda2
port 1175 nsew power bidirectional
rlabel metal5 s -8576 336676 592500 337276 6 vdda2
port 1176 nsew power bidirectional
rlabel metal5 s -8576 300676 592500 301276 6 vdda2
port 1177 nsew power bidirectional
rlabel metal5 s -8576 264676 592500 265276 6 vdda2
port 1178 nsew power bidirectional
rlabel metal5 s -8576 228676 592500 229276 6 vdda2
port 1179 nsew power bidirectional
rlabel metal5 s -8576 192676 592500 193276 6 vdda2
port 1180 nsew power bidirectional
rlabel metal5 s -8576 156676 592500 157276 6 vdda2
port 1181 nsew power bidirectional
rlabel metal5 s -8576 120676 592500 121276 6 vdda2
port 1182 nsew power bidirectional
rlabel metal5 s -8576 84676 592500 85276 6 vdda2
port 1183 nsew power bidirectional
rlabel metal5 s -8576 48676 592500 49276 6 vdda2
port 1184 nsew power bidirectional
rlabel metal5 s -8576 12676 592500 13276 6 vdda2
port 1185 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 1186 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 1187 nsew ground bidirectional
rlabel metal4 s 569604 693500 570204 711440 6 vssa2
port 1188 nsew ground bidirectional
rlabel metal4 s 533604 693500 534204 711440 6 vssa2
port 1189 nsew ground bidirectional
rlabel metal4 s 497604 693500 498204 711440 6 vssa2
port 1190 nsew ground bidirectional
rlabel metal4 s 461604 693500 462204 711440 6 vssa2
port 1191 nsew ground bidirectional
rlabel metal4 s 425604 693500 426204 711440 6 vssa2
port 1192 nsew ground bidirectional
rlabel metal4 s 389604 693500 390204 711440 6 vssa2
port 1193 nsew ground bidirectional
rlabel metal4 s 353604 693500 354204 711440 6 vssa2
port 1194 nsew ground bidirectional
rlabel metal4 s 317604 693500 318204 711440 6 vssa2
port 1195 nsew ground bidirectional
rlabel metal4 s 281604 693500 282204 711440 6 vssa2
port 1196 nsew ground bidirectional
rlabel metal4 s 245604 693500 246204 711440 6 vssa2
port 1197 nsew ground bidirectional
rlabel metal4 s 209604 693500 210204 711440 6 vssa2
port 1198 nsew ground bidirectional
rlabel metal4 s 173604 693500 174204 711440 6 vssa2
port 1199 nsew ground bidirectional
rlabel metal4 s 137604 693500 138204 711440 6 vssa2
port 1200 nsew ground bidirectional
rlabel metal4 s 101604 693500 102204 711440 6 vssa2
port 1201 nsew ground bidirectional
rlabel metal4 s 65604 693500 66204 711440 6 vssa2
port 1202 nsew ground bidirectional
rlabel metal4 s 29604 693500 30204 711440 6 vssa2
port 1203 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 1204 nsew ground bidirectional
rlabel metal4 s 569604 503500 570204 534500 6 vssa2
port 1205 nsew ground bidirectional
rlabel metal4 s 533604 503500 534204 534500 6 vssa2
port 1206 nsew ground bidirectional
rlabel metal4 s 497604 503500 498204 534500 6 vssa2
port 1207 nsew ground bidirectional
rlabel metal4 s 461604 503500 462204 534500 6 vssa2
port 1208 nsew ground bidirectional
rlabel metal4 s 425604 503500 426204 534500 6 vssa2
port 1209 nsew ground bidirectional
rlabel metal4 s 389604 249500 390204 534500 6 vssa2
port 1210 nsew ground bidirectional
rlabel metal4 s 353604 249500 354204 534500 6 vssa2
port 1211 nsew ground bidirectional
rlabel metal4 s 317604 -7504 318204 534500 6 vssa2
port 1212 nsew ground bidirectional
rlabel metal4 s 281604 -7504 282204 534500 6 vssa2
port 1213 nsew ground bidirectional
rlabel metal4 s 245604 -7504 246204 534500 6 vssa2
port 1214 nsew ground bidirectional
rlabel metal4 s 209604 249500 210204 534500 6 vssa2
port 1215 nsew ground bidirectional
rlabel metal4 s 173604 249500 174204 534500 6 vssa2
port 1216 nsew ground bidirectional
rlabel metal4 s 137604 493500 138204 534500 6 vssa2
port 1217 nsew ground bidirectional
rlabel metal4 s 101604 493500 102204 534500 6 vssa2
port 1218 nsew ground bidirectional
rlabel metal4 s 65604 493500 66204 534500 6 vssa2
port 1219 nsew ground bidirectional
rlabel metal4 s 29604 493500 30204 534500 6 vssa2
port 1220 nsew ground bidirectional
rlabel metal4 s 137604 249500 138204 338500 6 vssa2
port 1221 nsew ground bidirectional
rlabel metal4 s 101604 249500 102204 338500 6 vssa2
port 1222 nsew ground bidirectional
rlabel metal4 s 65604 249500 66204 338500 6 vssa2
port 1223 nsew ground bidirectional
rlabel metal4 s 29604 249500 30204 338500 6 vssa2
port 1224 nsew ground bidirectional
rlabel metal4 s 569604 249500 570204 334500 6 vssa2
port 1225 nsew ground bidirectional
rlabel metal4 s 533604 249500 534204 334500 6 vssa2
port 1226 nsew ground bidirectional
rlabel metal4 s 497604 249500 498204 334500 6 vssa2
port 1227 nsew ground bidirectional
rlabel metal4 s 461604 249500 462204 334500 6 vssa2
port 1228 nsew ground bidirectional
rlabel metal4 s 425604 249500 426204 334500 6 vssa2
port 1229 nsew ground bidirectional
rlabel metal4 s 569604 -7504 570204 10500 6 vssa2
port 1230 nsew ground bidirectional
rlabel metal4 s 533604 -7504 534204 10500 6 vssa2
port 1231 nsew ground bidirectional
rlabel metal4 s 497604 -7504 498204 10500 6 vssa2
port 1232 nsew ground bidirectional
rlabel metal4 s 461604 -7504 462204 10500 6 vssa2
port 1233 nsew ground bidirectional
rlabel metal4 s 425604 -7504 426204 10500 6 vssa2
port 1234 nsew ground bidirectional
rlabel metal4 s 389604 -7504 390204 10500 6 vssa2
port 1235 nsew ground bidirectional
rlabel metal4 s 353604 -7504 354204 10500 6 vssa2
port 1236 nsew ground bidirectional
rlabel metal4 s 209604 -7504 210204 10500 6 vssa2
port 1237 nsew ground bidirectional
rlabel metal4 s 173604 -7504 174204 10500 6 vssa2
port 1238 nsew ground bidirectional
rlabel metal4 s 137604 -7504 138204 10500 6 vssa2
port 1239 nsew ground bidirectional
rlabel metal4 s 101604 -7504 102204 10500 6 vssa2
port 1240 nsew ground bidirectional
rlabel metal4 s 65604 -7504 66204 10500 6 vssa2
port 1241 nsew ground bidirectional
rlabel metal4 s 29604 -7504 30204 10500 6 vssa2
port 1242 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 1243 nsew ground bidirectional
rlabel metal5 s -8576 678676 592500 679276 6 vssa2
port 1244 nsew ground bidirectional
rlabel metal5 s -8576 642676 592500 643276 6 vssa2
port 1245 nsew ground bidirectional
rlabel metal5 s -8576 606676 592500 607276 6 vssa2
port 1246 nsew ground bidirectional
rlabel metal5 s -8576 570676 592500 571276 6 vssa2
port 1247 nsew ground bidirectional
rlabel metal5 s -8576 534676 592500 535276 6 vssa2
port 1248 nsew ground bidirectional
rlabel metal5 s -8576 498676 592500 499276 6 vssa2
port 1249 nsew ground bidirectional
rlabel metal5 s -8576 462676 592500 463276 6 vssa2
port 1250 nsew ground bidirectional
rlabel metal5 s -8576 426676 592500 427276 6 vssa2
port 1251 nsew ground bidirectional
rlabel metal5 s -8576 390676 592500 391276 6 vssa2
port 1252 nsew ground bidirectional
rlabel metal5 s -8576 354676 592500 355276 6 vssa2
port 1253 nsew ground bidirectional
rlabel metal5 s -8576 318676 592500 319276 6 vssa2
port 1254 nsew ground bidirectional
rlabel metal5 s -8576 282676 592500 283276 6 vssa2
port 1255 nsew ground bidirectional
rlabel metal5 s -8576 246676 592500 247276 6 vssa2
port 1256 nsew ground bidirectional
rlabel metal5 s -8576 210676 592500 211276 6 vssa2
port 1257 nsew ground bidirectional
rlabel metal5 s -8576 174676 592500 175276 6 vssa2
port 1258 nsew ground bidirectional
rlabel metal5 s -8576 138676 592500 139276 6 vssa2
port 1259 nsew ground bidirectional
rlabel metal5 s -8576 102676 592500 103276 6 vssa2
port 1260 nsew ground bidirectional
rlabel metal5 s -8576 66676 592500 67276 6 vssa2
port 1261 nsew ground bidirectional
rlabel metal5 s -8576 30676 592500 31276 6 vssa2
port 1262 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 1263 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 584000 704000
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 908860280
string GDS_START 723796886
<< end >>

