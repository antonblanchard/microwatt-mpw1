VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_512x64
  CLASS BLOCK ;
  FOREIGN RAM_512x64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 700.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2447.290 0.000 2447.570 4.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.150 0.000 2466.430 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.470 0.000 2485.750 4.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2504.330 0.000 2504.610 4.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2523.190 0.000 2523.470 4.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2542.510 0.000 2542.790 4.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2561.370 0.000 2561.650 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2580.690 0.000 2580.970 4.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2599.550 0.000 2599.830 4.000 ;
    END
  END A[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2618.410 0.000 2618.690 4.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.290 0.000 1228.570 4.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 0.000 1419.010 4.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.590 0.000 1437.870 4.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.910 0.000 1457.190 4.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.770 0.000 1476.050 4.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.630 0.000 1494.910 4.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.950 0.000 1514.230 4.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 0.000 1533.090 4.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.990 0.000 1571.270 4.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.850 0.000 1590.130 4.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 4.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.170 0.000 1609.450 4.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.030 0.000 1628.310 4.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.350 0.000 1647.630 4.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.210 0.000 1666.490 4.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.070 0.000 1685.350 4.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.390 0.000 1704.670 4.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.250 0.000 1723.530 4.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.570 0.000 1742.850 4.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 0.000 1761.710 4.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.290 0.000 1780.570 4.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.610 0.000 1799.890 4.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.470 0.000 1818.750 4.000 ;
    END
  END Di[31]
  PIN Di[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.790 0.000 1838.070 4.000 ;
    END
  END Di[32]
  PIN Di[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1856.650 0.000 1856.930 4.000 ;
    END
  END Di[33]
  PIN Di[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.970 0.000 1876.250 4.000 ;
    END
  END Di[34]
  PIN Di[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.830 0.000 1895.110 4.000 ;
    END
  END Di[35]
  PIN Di[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.690 0.000 1913.970 4.000 ;
    END
  END Di[36]
  PIN Di[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.010 0.000 1933.290 4.000 ;
    END
  END Di[37]
  PIN Di[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.870 0.000 1952.150 4.000 ;
    END
  END Di[38]
  PIN Di[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.190 0.000 1971.470 4.000 ;
    END
  END Di[39]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.330 0.000 1285.610 4.000 ;
    END
  END Di[3]
  PIN Di[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.050 0.000 1990.330 4.000 ;
    END
  END Di[40]
  PIN Di[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.910 0.000 2009.190 4.000 ;
    END
  END Di[41]
  PIN Di[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.230 0.000 2028.510 4.000 ;
    END
  END Di[42]
  PIN Di[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.090 0.000 2047.370 4.000 ;
    END
  END Di[43]
  PIN Di[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.410 0.000 2066.690 4.000 ;
    END
  END Di[44]
  PIN Di[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.270 0.000 2085.550 4.000 ;
    END
  END Di[45]
  PIN Di[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2104.130 0.000 2104.410 4.000 ;
    END
  END Di[46]
  PIN Di[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2123.450 0.000 2123.730 4.000 ;
    END
  END Di[47]
  PIN Di[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.310 0.000 2142.590 4.000 ;
    END
  END Di[48]
  PIN Di[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.630 0.000 2161.910 4.000 ;
    END
  END Di[49]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 0.000 1304.470 4.000 ;
    END
  END Di[4]
  PIN Di[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.490 0.000 2180.770 4.000 ;
    END
  END Di[50]
  PIN Di[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.350 0.000 2199.630 4.000 ;
    END
  END Di[51]
  PIN Di[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.670 0.000 2218.950 4.000 ;
    END
  END Di[52]
  PIN Di[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.530 0.000 2237.810 4.000 ;
    END
  END Di[53]
  PIN Di[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.850 0.000 2257.130 4.000 ;
    END
  END Di[54]
  PIN Di[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2275.710 0.000 2275.990 4.000 ;
    END
  END Di[55]
  PIN Di[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2294.570 0.000 2294.850 4.000 ;
    END
  END Di[56]
  PIN Di[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.890 0.000 2314.170 4.000 ;
    END
  END Di[57]
  PIN Di[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2332.750 0.000 2333.030 4.000 ;
    END
  END Di[58]
  PIN Di[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2352.070 0.000 2352.350 4.000 ;
    END
  END Di[59]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END Di[5]
  PIN Di[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.930 0.000 2371.210 4.000 ;
    END
  END Di[60]
  PIN Di[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.250 0.000 2390.530 4.000 ;
    END
  END Di[61]
  PIN Di[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2409.110 0.000 2409.390 4.000 ;
    END
  END Di[62]
  PIN Di[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2427.970 0.000 2428.250 4.000 ;
    END
  END Di[63]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1361.230 0.000 1361.510 4.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.550 0.000 1380.830 4.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.410 0.000 1399.690 4.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END Do[31]
  PIN Do[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END Do[32]
  PIN Do[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END Do[33]
  PIN Do[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END Do[34]
  PIN Do[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 0.000 676.110 4.000 ;
    END
  END Do[35]
  PIN Do[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 0.000 694.970 4.000 ;
    END
  END Do[36]
  PIN Do[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END Do[37]
  PIN Do[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END Do[38]
  PIN Do[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 0.000 752.010 4.000 ;
    END
  END Do[39]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END Do[3]
  PIN Do[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END Do[40]
  PIN Do[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END Do[41]
  PIN Do[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 0.000 809.510 4.000 ;
    END
  END Do[42]
  PIN Do[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 4.000 ;
    END
  END Do[43]
  PIN Do[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END Do[44]
  PIN Do[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END Do[45]
  PIN Do[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 0.000 885.410 4.000 ;
    END
  END Do[46]
  PIN Do[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.450 0.000 904.730 4.000 ;
    END
  END Do[47]
  PIN Do[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.310 0.000 923.590 4.000 ;
    END
  END Do[48]
  PIN Do[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 0.000 942.910 4.000 ;
    END
  END Do[49]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END Do[4]
  PIN Do[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 0.000 961.770 4.000 ;
    END
  END Do[50]
  PIN Do[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END Do[51]
  PIN Do[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 4.000 ;
    END
  END Do[52]
  PIN Do[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.530 0.000 1018.810 4.000 ;
    END
  END Do[53]
  PIN Do[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 0.000 1038.130 4.000 ;
    END
  END Do[54]
  PIN Do[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 0.000 1056.990 4.000 ;
    END
  END Do[55]
  PIN Do[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END Do[56]
  PIN Do[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END Do[57]
  PIN Do[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.750 0.000 1114.030 4.000 ;
    END
  END Do[58]
  PIN Do[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.070 0.000 1133.350 4.000 ;
    END
  END Do[59]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END Do[5]
  PIN Do[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END Do[60]
  PIN Do[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.790 0.000 1171.070 4.000 ;
    END
  END Do[61]
  PIN Do[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.110 0.000 1190.390 4.000 ;
    END
  END Do[62]
  PIN Do[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 0.000 1209.250 4.000 ;
    END
  END Do[63]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2789.990 0.000 2790.270 4.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2637.730 0.000 2638.010 4.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.590 0.000 2656.870 4.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2675.910 0.000 2676.190 4.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2694.770 0.000 2695.050 4.000 ;
    END
  END WE[3]
  PIN WE[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2713.630 0.000 2713.910 4.000 ;
    END
  END WE[4]
  PIN WE[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.950 0.000 2733.230 4.000 ;
    END
  END WE[5]
  PIN WE[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.810 0.000 2752.090 4.000 ;
    END
  END WE[6]
  PIN WE[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2771.130 0.000 2771.410 4.000 ;
    END
  END WE[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 686.805 1047.955 686.855 ;
        RECT 5.330 684.075 2794.230 686.805 ;
        RECT 5.330 684.025 660.635 684.075 ;
        RECT 5.330 681.365 93.455 681.415 ;
        RECT 5.330 678.635 2794.230 681.365 ;
        RECT 5.330 678.585 175.335 678.635 ;
        RECT 5.330 675.925 120.595 675.975 ;
        RECT 5.330 673.195 2794.230 675.925 ;
        RECT 5.330 673.145 56.195 673.195 ;
        RECT 5.330 670.485 248.935 670.535 ;
        RECT 5.330 667.755 2794.230 670.485 ;
        RECT 5.330 667.705 147.275 667.755 ;
        RECT 5.330 665.045 165.215 665.095 ;
        RECT 5.330 662.315 2794.230 665.045 ;
        RECT 5.330 662.265 137.155 662.315 ;
        RECT 5.330 659.605 640.855 659.655 ;
        RECT 5.330 656.875 2794.230 659.605 ;
        RECT 5.330 656.825 180.395 656.875 ;
        RECT 5.330 654.165 715.375 654.215 ;
        RECT 5.330 651.435 2794.230 654.165 ;
        RECT 5.330 651.385 203.395 651.435 ;
        RECT 5.330 648.725 374.515 648.775 ;
        RECT 5.330 645.995 2794.230 648.725 ;
        RECT 5.330 645.945 119.215 645.995 ;
        RECT 5.330 643.285 536.895 643.335 ;
        RECT 5.330 640.555 2794.230 643.285 ;
        RECT 5.330 640.505 345.075 640.555 ;
        RECT 5.330 637.845 470.195 637.895 ;
        RECT 5.330 635.115 2794.230 637.845 ;
        RECT 5.330 635.065 119.215 635.115 ;
        RECT 5.330 632.405 230.075 632.455 ;
        RECT 5.330 629.675 2794.230 632.405 ;
        RECT 5.330 629.625 190.515 629.675 ;
        RECT 5.330 626.965 174.415 627.015 ;
        RECT 5.330 624.235 2794.230 626.965 ;
        RECT 5.330 624.185 181.315 624.235 ;
        RECT 5.330 621.525 84.715 621.575 ;
        RECT 5.330 618.795 2794.230 621.525 ;
        RECT 5.330 618.745 251.695 618.795 ;
        RECT 5.330 616.085 77.355 616.135 ;
        RECT 5.330 613.355 2794.230 616.085 ;
        RECT 5.330 613.305 165.675 613.355 ;
        RECT 5.330 610.645 105.415 610.695 ;
        RECT 5.330 607.915 2794.230 610.645 ;
        RECT 5.330 607.865 231.455 607.915 ;
        RECT 5.330 605.205 105.415 605.255 ;
        RECT 5.330 602.475 2794.230 605.205 ;
        RECT 5.330 602.425 222.255 602.475 ;
        RECT 5.330 599.765 200.635 599.815 ;
        RECT 5.330 597.035 2794.230 599.765 ;
        RECT 5.330 596.985 188.675 597.035 ;
        RECT 5.330 594.325 60.795 594.375 ;
        RECT 5.330 591.595 2794.230 594.325 ;
        RECT 5.330 591.545 84.255 591.595 ;
        RECT 5.330 588.885 222.715 588.935 ;
        RECT 5.330 586.155 2794.230 588.885 ;
        RECT 5.330 586.105 287.575 586.155 ;
        RECT 5.330 583.445 178.555 583.495 ;
        RECT 5.330 580.715 2794.230 583.445 ;
        RECT 5.330 580.665 41.015 580.715 ;
        RECT 5.330 578.005 105.415 578.055 ;
        RECT 5.330 575.275 2794.230 578.005 ;
        RECT 5.330 575.225 147.275 575.275 ;
        RECT 5.330 572.565 126.575 572.615 ;
        RECT 5.330 569.835 2794.230 572.565 ;
        RECT 5.330 569.785 126.115 569.835 ;
        RECT 5.330 567.125 210.755 567.175 ;
        RECT 5.330 564.395 2794.230 567.125 ;
        RECT 5.330 564.345 165.215 564.395 ;
        RECT 5.330 561.685 306.435 561.735 ;
        RECT 5.330 558.955 2794.230 561.685 ;
        RECT 5.330 558.905 119.215 558.955 ;
        RECT 5.330 556.245 91.155 556.295 ;
        RECT 5.330 553.515 2794.230 556.245 ;
        RECT 5.330 553.465 361.635 553.515 ;
        RECT 5.330 550.805 218.575 550.855 ;
        RECT 5.330 548.075 2794.230 550.805 ;
        RECT 5.330 548.025 140.375 548.075 ;
        RECT 5.330 545.365 423.735 545.415 ;
        RECT 5.330 542.635 2794.230 545.365 ;
        RECT 5.330 542.585 124.735 542.635 ;
        RECT 5.330 539.925 294.015 539.975 ;
        RECT 5.330 537.195 2794.230 539.925 ;
        RECT 5.330 537.145 111.855 537.195 ;
        RECT 5.330 534.485 501.935 534.535 ;
        RECT 5.330 531.755 2794.230 534.485 ;
        RECT 5.330 531.705 101.275 531.755 ;
        RECT 5.330 529.045 225.475 529.095 ;
        RECT 5.330 526.315 2794.230 529.045 ;
        RECT 5.330 526.265 441.675 526.315 ;
        RECT 5.330 523.605 77.355 523.655 ;
        RECT 5.330 520.875 2794.230 523.605 ;
        RECT 5.330 520.825 189.135 520.875 ;
        RECT 5.330 518.165 108.175 518.215 ;
        RECT 5.330 515.435 2794.230 518.165 ;
        RECT 5.330 515.385 147.275 515.435 ;
        RECT 5.330 512.725 204.315 512.775 ;
        RECT 5.330 509.995 2794.230 512.725 ;
        RECT 5.330 509.945 149.575 509.995 ;
        RECT 5.330 507.285 113.235 507.335 ;
        RECT 5.330 504.555 2794.230 507.285 ;
        RECT 5.330 504.505 317.015 504.555 ;
        RECT 5.330 501.845 414.075 501.895 ;
        RECT 5.330 499.115 2794.230 501.845 ;
        RECT 5.330 499.065 224.555 499.115 ;
        RECT 5.330 496.405 245.715 496.455 ;
        RECT 5.330 493.675 2794.230 496.405 ;
        RECT 5.330 493.625 371.755 493.675 ;
        RECT 5.330 490.965 114.615 491.015 ;
        RECT 5.330 488.235 2794.230 490.965 ;
        RECT 5.330 488.185 92.995 488.235 ;
        RECT 5.330 485.525 84.715 485.575 ;
        RECT 5.330 482.795 2794.230 485.525 ;
        RECT 5.330 482.745 483.995 482.795 ;
        RECT 5.330 480.085 230.075 480.135 ;
        RECT 5.330 477.355 2794.230 480.085 ;
        RECT 5.330 477.305 136.235 477.355 ;
        RECT 5.330 474.645 173.495 474.695 ;
        RECT 5.330 471.915 2794.230 474.645 ;
        RECT 5.330 471.865 81.495 471.915 ;
        RECT 5.330 469.205 161.535 469.255 ;
        RECT 5.330 466.475 2794.230 469.205 ;
        RECT 5.330 466.425 179.475 466.475 ;
        RECT 5.330 463.765 107.715 463.815 ;
        RECT 5.330 461.035 2794.230 463.765 ;
        RECT 5.330 460.985 512.055 461.035 ;
        RECT 5.330 458.325 470.195 458.375 ;
        RECT 5.330 455.595 2794.230 458.325 ;
        RECT 5.330 455.545 91.155 455.595 ;
        RECT 5.330 452.885 121.975 452.935 ;
        RECT 5.330 450.155 2794.230 452.885 ;
        RECT 5.330 450.105 97.135 450.155 ;
        RECT 5.330 447.445 121.975 447.495 ;
        RECT 5.330 444.715 2794.230 447.445 ;
        RECT 5.330 444.665 262.735 444.715 ;
        RECT 5.330 442.005 57.115 442.055 ;
        RECT 5.330 439.275 2794.230 442.005 ;
        RECT 5.330 439.225 102.655 439.275 ;
        RECT 5.330 436.565 92.995 436.615 ;
        RECT 5.330 433.835 2794.230 436.565 ;
        RECT 5.330 433.785 360.255 433.835 ;
        RECT 5.330 431.125 126.575 431.175 ;
        RECT 5.330 428.395 2794.230 431.125 ;
        RECT 5.330 428.345 91.155 428.395 ;
        RECT 5.330 425.685 126.575 425.735 ;
        RECT 5.330 422.955 2794.230 425.685 ;
        RECT 5.330 422.905 70.455 422.955 ;
        RECT 5.330 420.245 95.295 420.295 ;
        RECT 5.330 417.515 2794.230 420.245 ;
        RECT 5.330 417.465 105.415 417.515 ;
        RECT 5.330 414.805 121.515 414.855 ;
        RECT 5.330 412.075 2794.230 414.805 ;
        RECT 5.330 412.025 299.995 412.075 ;
        RECT 5.330 409.365 64.475 409.415 ;
        RECT 5.330 406.635 2794.230 409.365 ;
        RECT 5.330 406.585 76.895 406.635 ;
        RECT 5.330 403.925 94.835 403.975 ;
        RECT 5.330 401.195 2794.230 403.925 ;
        RECT 5.330 401.145 131.635 401.195 ;
        RECT 5.330 398.485 217.655 398.535 ;
        RECT 5.330 395.755 2794.230 398.485 ;
        RECT 5.330 395.705 316.555 395.755 ;
        RECT 5.330 393.045 491.355 393.095 ;
        RECT 5.330 390.315 2794.230 393.045 ;
        RECT 5.330 390.265 491.815 390.315 ;
        RECT 5.330 387.605 995.515 387.655 ;
        RECT 5.330 384.875 2794.230 387.605 ;
        RECT 5.330 384.825 828.535 384.875 ;
        RECT 5.330 382.165 77.355 382.215 ;
        RECT 5.330 379.435 2794.230 382.165 ;
        RECT 5.330 379.385 166.595 379.435 ;
        RECT 5.330 376.725 93.455 376.775 ;
        RECT 5.330 373.995 2794.230 376.725 ;
        RECT 5.330 373.945 98.515 373.995 ;
        RECT 5.330 371.285 62.175 371.335 ;
        RECT 5.330 368.555 2794.230 371.285 ;
        RECT 5.330 368.505 35.495 368.555 ;
        RECT 5.330 365.845 596.695 365.895 ;
        RECT 5.330 363.115 2794.230 365.845 ;
        RECT 5.330 363.065 148.195 363.115 ;
        RECT 5.330 360.405 105.415 360.455 ;
        RECT 5.330 357.675 2794.230 360.405 ;
        RECT 5.330 357.625 103.575 357.675 ;
        RECT 5.330 354.965 143.135 355.015 ;
        RECT 5.330 352.235 2794.230 354.965 ;
        RECT 5.330 352.185 63.095 352.235 ;
        RECT 5.330 349.525 84.715 349.575 ;
        RECT 5.330 346.795 2794.230 349.525 ;
        RECT 5.330 346.745 111.395 346.795 ;
        RECT 5.330 344.085 105.415 344.135 ;
        RECT 5.330 341.355 2794.230 344.085 ;
        RECT 5.330 341.305 403.495 341.355 ;
        RECT 5.330 338.645 81.955 338.695 ;
        RECT 5.330 335.915 2794.230 338.645 ;
        RECT 5.330 335.865 149.575 335.915 ;
        RECT 5.330 333.205 115.535 333.255 ;
        RECT 5.330 330.475 2794.230 333.205 ;
        RECT 5.330 330.425 56.195 330.475 ;
        RECT 5.330 327.765 144.515 327.815 ;
        RECT 5.330 325.035 2794.230 327.765 ;
        RECT 5.330 324.985 147.275 325.035 ;
        RECT 5.330 322.325 35.035 322.375 ;
        RECT 5.330 319.595 2794.230 322.325 ;
        RECT 5.330 319.545 119.215 319.595 ;
        RECT 5.330 316.885 144.975 316.935 ;
        RECT 5.330 314.155 2794.230 316.885 ;
        RECT 5.330 314.105 108.635 314.155 ;
        RECT 5.330 311.445 121.055 311.495 ;
        RECT 5.330 308.715 2794.230 311.445 ;
        RECT 5.330 308.665 12.035 308.715 ;
        RECT 5.330 306.005 1148.695 306.055 ;
        RECT 5.330 303.275 2794.230 306.005 ;
        RECT 5.330 303.225 588.875 303.275 ;
        RECT 5.330 300.565 489.515 300.615 ;
        RECT 5.330 297.835 2794.230 300.565 ;
        RECT 5.330 297.785 64.015 297.835 ;
        RECT 5.330 295.125 181.775 295.175 ;
        RECT 5.330 292.395 2794.230 295.125 ;
        RECT 5.330 292.345 16.635 292.395 ;
        RECT 5.330 289.685 229.615 289.735 ;
        RECT 5.330 286.955 2794.230 289.685 ;
        RECT 5.330 286.905 409.935 286.955 ;
        RECT 5.330 284.245 120.595 284.295 ;
        RECT 5.330 281.515 2794.230 284.245 ;
        RECT 5.330 281.465 79.195 281.515 ;
        RECT 5.330 278.805 105.415 278.855 ;
        RECT 5.330 276.075 2794.230 278.805 ;
        RECT 5.330 276.025 64.015 276.075 ;
        RECT 5.330 273.365 113.695 273.415 ;
        RECT 5.330 270.635 2794.230 273.365 ;
        RECT 5.330 270.585 298.155 270.635 ;
        RECT 5.330 267.925 133.475 267.975 ;
        RECT 5.330 265.195 2794.230 267.925 ;
        RECT 5.330 265.145 196.495 265.195 ;
        RECT 5.330 262.485 115.075 262.535 ;
        RECT 5.330 259.755 2794.230 262.485 ;
        RECT 5.330 259.705 203.395 259.755 ;
        RECT 5.330 257.045 135.775 257.095 ;
        RECT 5.330 254.315 2794.230 257.045 ;
        RECT 5.330 254.265 122.895 254.315 ;
        RECT 5.330 251.605 68.615 251.655 ;
        RECT 5.330 248.875 2794.230 251.605 ;
        RECT 5.330 248.825 74.135 248.875 ;
        RECT 5.330 246.165 62.635 246.215 ;
        RECT 5.330 243.435 2794.230 246.165 ;
        RECT 5.330 243.385 119.215 243.435 ;
        RECT 5.330 240.725 49.755 240.775 ;
        RECT 5.330 237.995 2794.230 240.725 ;
        RECT 5.330 237.945 51.135 237.995 ;
        RECT 5.330 235.285 919.155 235.335 ;
        RECT 5.330 232.555 2794.230 235.285 ;
        RECT 5.330 232.505 215.815 232.555 ;
        RECT 5.330 229.845 345.995 229.895 ;
        RECT 5.330 227.115 2794.230 229.845 ;
        RECT 5.330 227.065 165.215 227.115 ;
        RECT 5.330 224.405 112.775 224.455 ;
        RECT 5.330 221.675 2794.230 224.405 ;
        RECT 5.330 221.625 98.975 221.675 ;
        RECT 5.330 218.965 94.375 219.015 ;
        RECT 5.330 216.235 2794.230 218.965 ;
        RECT 5.330 216.185 119.215 216.235 ;
        RECT 5.330 213.525 562.655 213.575 ;
        RECT 5.330 210.795 2794.230 213.525 ;
        RECT 5.330 210.745 353.355 210.795 ;
        RECT 5.330 208.085 85.175 208.135 ;
        RECT 5.330 205.355 2794.230 208.085 ;
        RECT 5.330 205.305 94.375 205.355 ;
        RECT 5.330 202.645 219.035 202.695 ;
        RECT 5.330 199.915 2794.230 202.645 ;
        RECT 5.330 199.865 52.055 199.915 ;
        RECT 5.330 197.205 126.115 197.255 ;
        RECT 5.330 194.475 2794.230 197.205 ;
        RECT 5.330 194.425 97.595 194.475 ;
        RECT 5.330 191.765 95.755 191.815 ;
        RECT 5.330 189.035 2794.230 191.765 ;
        RECT 5.330 188.985 359.335 189.035 ;
        RECT 5.330 186.325 217.655 186.375 ;
        RECT 5.330 183.595 2794.230 186.325 ;
        RECT 5.330 183.545 391.535 183.595 ;
        RECT 5.330 180.885 391.535 180.935 ;
        RECT 5.330 178.155 2794.230 180.885 ;
        RECT 5.330 178.105 136.695 178.155 ;
        RECT 5.330 175.445 42.395 175.495 ;
        RECT 5.330 172.715 2794.230 175.445 ;
        RECT 5.330 172.665 427.875 172.715 ;
        RECT 5.330 170.005 245.715 170.055 ;
        RECT 5.330 167.275 2794.230 170.005 ;
        RECT 5.330 167.225 157.855 167.275 ;
        RECT 5.330 164.565 233.755 164.615 ;
        RECT 5.330 161.835 2794.230 164.565 ;
        RECT 5.330 161.785 41.015 161.835 ;
        RECT 5.330 159.125 217.655 159.175 ;
        RECT 5.330 156.395 2794.230 159.125 ;
        RECT 5.330 156.345 63.095 156.395 ;
        RECT 5.330 153.685 194.655 153.735 ;
        RECT 5.330 150.955 2794.230 153.685 ;
        RECT 5.330 150.905 108.635 150.955 ;
        RECT 5.330 148.245 140.835 148.295 ;
        RECT 5.330 145.515 2794.230 148.245 ;
        RECT 5.330 145.465 35.035 145.515 ;
        RECT 5.330 142.805 373.595 142.855 ;
        RECT 5.330 140.075 2794.230 142.805 ;
        RECT 5.330 140.025 110.015 140.075 ;
        RECT 5.330 137.365 124.275 137.415 ;
        RECT 5.330 134.635 2794.230 137.365 ;
        RECT 5.330 134.585 119.215 134.635 ;
        RECT 5.330 131.925 66.775 131.975 ;
        RECT 5.330 129.195 2794.230 131.925 ;
        RECT 5.330 129.145 175.335 129.195 ;
        RECT 5.330 126.485 193.275 126.535 ;
        RECT 5.330 123.755 2794.230 126.485 ;
        RECT 5.330 123.705 203.395 123.755 ;
        RECT 5.330 121.045 49.295 121.095 ;
        RECT 5.330 118.315 2794.230 121.045 ;
        RECT 5.330 118.265 91.155 118.315 ;
        RECT 5.330 115.605 86.555 115.655 ;
        RECT 5.330 112.875 2794.230 115.605 ;
        RECT 5.330 112.825 210.755 112.875 ;
        RECT 5.330 110.165 105.415 110.215 ;
        RECT 5.330 107.435 2794.230 110.165 ;
        RECT 5.330 107.385 44.235 107.435 ;
        RECT 5.330 104.725 161.535 104.775 ;
        RECT 5.330 101.995 2794.230 104.725 ;
        RECT 5.330 101.945 137.615 101.995 ;
        RECT 5.330 99.285 199.715 99.335 ;
        RECT 5.330 96.555 2794.230 99.285 ;
        RECT 5.330 96.505 147.275 96.555 ;
        RECT 5.330 93.845 424.655 93.895 ;
        RECT 5.330 91.115 2794.230 93.845 ;
        RECT 5.330 91.065 315.635 91.115 ;
        RECT 5.330 88.405 57.575 88.455 ;
        RECT 5.330 85.675 2794.230 88.405 ;
        RECT 5.330 85.625 91.155 85.675 ;
        RECT 5.330 82.965 31.815 83.015 ;
        RECT 5.330 80.235 2794.230 82.965 ;
        RECT 5.330 80.185 308.735 80.235 ;
        RECT 5.330 77.525 136.235 77.575 ;
        RECT 5.330 74.795 2794.230 77.525 ;
        RECT 5.330 74.745 48.375 74.795 ;
        RECT 5.330 72.085 113.695 72.135 ;
        RECT 5.330 69.355 2794.230 72.085 ;
        RECT 5.330 69.305 119.215 69.355 ;
        RECT 5.330 66.645 38.715 66.695 ;
        RECT 5.330 63.915 2794.230 66.645 ;
        RECT 5.330 63.865 203.395 63.915 ;
        RECT 5.330 61.205 140.835 61.255 ;
        RECT 5.330 58.475 2794.230 61.205 ;
        RECT 5.330 58.425 43.315 58.475 ;
        RECT 5.330 55.765 311.495 55.815 ;
        RECT 5.330 53.035 2794.230 55.765 ;
        RECT 5.330 52.985 12.955 53.035 ;
        RECT 5.330 50.325 189.595 50.375 ;
        RECT 5.330 47.595 2794.230 50.325 ;
        RECT 5.330 47.545 49.295 47.595 ;
        RECT 5.330 44.885 92.075 44.935 ;
        RECT 5.330 42.155 2794.230 44.885 ;
        RECT 5.330 42.105 128.875 42.155 ;
        RECT 5.330 39.445 115.535 39.495 ;
        RECT 5.330 36.715 2794.230 39.445 ;
        RECT 5.330 36.665 100.355 36.715 ;
        RECT 5.330 34.005 225.015 34.055 ;
        RECT 5.330 31.275 2794.230 34.005 ;
        RECT 5.330 31.225 241.575 31.275 ;
        RECT 5.330 28.565 340.475 28.615 ;
        RECT 5.330 25.835 2794.230 28.565 ;
        RECT 5.330 25.785 277.455 25.835 ;
        RECT 5.330 23.125 571.855 23.175 ;
        RECT 5.330 20.395 2794.230 23.125 ;
        RECT 5.330 20.345 820.715 20.395 ;
        RECT 5.330 17.685 1739.335 17.735 ;
        RECT 5.330 14.955 2794.230 17.685 ;
        RECT 5.330 14.905 950.895 14.955 ;
        RECT 5.330 10.690 2794.230 12.295 ;
      LAYER li1 ;
        RECT 5.520 6.545 2794.040 690.455 ;
      LAYER met1 ;
        RECT 5.520 5.820 2794.040 690.500 ;
      LAYER met2 ;
        RECT 9.300 4.280 2791.180 690.530 ;
        RECT 9.850 4.000 27.870 4.280 ;
        RECT 28.710 4.000 46.730 4.280 ;
        RECT 47.570 4.000 66.050 4.280 ;
        RECT 66.890 4.000 84.910 4.280 ;
        RECT 85.750 4.000 104.230 4.280 ;
        RECT 105.070 4.000 123.090 4.280 ;
        RECT 123.930 4.000 141.950 4.280 ;
        RECT 142.790 4.000 161.270 4.280 ;
        RECT 162.110 4.000 180.130 4.280 ;
        RECT 180.970 4.000 199.450 4.280 ;
        RECT 200.290 4.000 218.310 4.280 ;
        RECT 219.150 4.000 237.170 4.280 ;
        RECT 238.010 4.000 256.490 4.280 ;
        RECT 257.330 4.000 275.350 4.280 ;
        RECT 276.190 4.000 294.670 4.280 ;
        RECT 295.510 4.000 313.530 4.280 ;
        RECT 314.370 4.000 332.390 4.280 ;
        RECT 333.230 4.000 351.710 4.280 ;
        RECT 352.550 4.000 370.570 4.280 ;
        RECT 371.410 4.000 389.890 4.280 ;
        RECT 390.730 4.000 408.750 4.280 ;
        RECT 409.590 4.000 427.610 4.280 ;
        RECT 428.450 4.000 446.930 4.280 ;
        RECT 447.770 4.000 465.790 4.280 ;
        RECT 466.630 4.000 485.110 4.280 ;
        RECT 485.950 4.000 503.970 4.280 ;
        RECT 504.810 4.000 523.290 4.280 ;
        RECT 524.130 4.000 542.150 4.280 ;
        RECT 542.990 4.000 561.010 4.280 ;
        RECT 561.850 4.000 580.330 4.280 ;
        RECT 581.170 4.000 599.190 4.280 ;
        RECT 600.030 4.000 618.510 4.280 ;
        RECT 619.350 4.000 637.370 4.280 ;
        RECT 638.210 4.000 656.230 4.280 ;
        RECT 657.070 4.000 675.550 4.280 ;
        RECT 676.390 4.000 694.410 4.280 ;
        RECT 695.250 4.000 713.730 4.280 ;
        RECT 714.570 4.000 732.590 4.280 ;
        RECT 733.430 4.000 751.450 4.280 ;
        RECT 752.290 4.000 770.770 4.280 ;
        RECT 771.610 4.000 789.630 4.280 ;
        RECT 790.470 4.000 808.950 4.280 ;
        RECT 809.790 4.000 827.810 4.280 ;
        RECT 828.650 4.000 846.670 4.280 ;
        RECT 847.510 4.000 865.990 4.280 ;
        RECT 866.830 4.000 884.850 4.280 ;
        RECT 885.690 4.000 904.170 4.280 ;
        RECT 905.010 4.000 923.030 4.280 ;
        RECT 923.870 4.000 942.350 4.280 ;
        RECT 943.190 4.000 961.210 4.280 ;
        RECT 962.050 4.000 980.070 4.280 ;
        RECT 980.910 4.000 999.390 4.280 ;
        RECT 1000.230 4.000 1018.250 4.280 ;
        RECT 1019.090 4.000 1037.570 4.280 ;
        RECT 1038.410 4.000 1056.430 4.280 ;
        RECT 1057.270 4.000 1075.290 4.280 ;
        RECT 1076.130 4.000 1094.610 4.280 ;
        RECT 1095.450 4.000 1113.470 4.280 ;
        RECT 1114.310 4.000 1132.790 4.280 ;
        RECT 1133.630 4.000 1151.650 4.280 ;
        RECT 1152.490 4.000 1170.510 4.280 ;
        RECT 1171.350 4.000 1189.830 4.280 ;
        RECT 1190.670 4.000 1208.690 4.280 ;
        RECT 1209.530 4.000 1228.010 4.280 ;
        RECT 1228.850 4.000 1246.870 4.280 ;
        RECT 1247.710 4.000 1265.730 4.280 ;
        RECT 1266.570 4.000 1285.050 4.280 ;
        RECT 1285.890 4.000 1303.910 4.280 ;
        RECT 1304.750 4.000 1323.230 4.280 ;
        RECT 1324.070 4.000 1342.090 4.280 ;
        RECT 1342.930 4.000 1360.950 4.280 ;
        RECT 1361.790 4.000 1380.270 4.280 ;
        RECT 1381.110 4.000 1399.130 4.280 ;
        RECT 1399.970 4.000 1418.450 4.280 ;
        RECT 1419.290 4.000 1437.310 4.280 ;
        RECT 1438.150 4.000 1456.630 4.280 ;
        RECT 1457.470 4.000 1475.490 4.280 ;
        RECT 1476.330 4.000 1494.350 4.280 ;
        RECT 1495.190 4.000 1513.670 4.280 ;
        RECT 1514.510 4.000 1532.530 4.280 ;
        RECT 1533.370 4.000 1551.850 4.280 ;
        RECT 1552.690 4.000 1570.710 4.280 ;
        RECT 1571.550 4.000 1589.570 4.280 ;
        RECT 1590.410 4.000 1608.890 4.280 ;
        RECT 1609.730 4.000 1627.750 4.280 ;
        RECT 1628.590 4.000 1647.070 4.280 ;
        RECT 1647.910 4.000 1665.930 4.280 ;
        RECT 1666.770 4.000 1684.790 4.280 ;
        RECT 1685.630 4.000 1704.110 4.280 ;
        RECT 1704.950 4.000 1722.970 4.280 ;
        RECT 1723.810 4.000 1742.290 4.280 ;
        RECT 1743.130 4.000 1761.150 4.280 ;
        RECT 1761.990 4.000 1780.010 4.280 ;
        RECT 1780.850 4.000 1799.330 4.280 ;
        RECT 1800.170 4.000 1818.190 4.280 ;
        RECT 1819.030 4.000 1837.510 4.280 ;
        RECT 1838.350 4.000 1856.370 4.280 ;
        RECT 1857.210 4.000 1875.690 4.280 ;
        RECT 1876.530 4.000 1894.550 4.280 ;
        RECT 1895.390 4.000 1913.410 4.280 ;
        RECT 1914.250 4.000 1932.730 4.280 ;
        RECT 1933.570 4.000 1951.590 4.280 ;
        RECT 1952.430 4.000 1970.910 4.280 ;
        RECT 1971.750 4.000 1989.770 4.280 ;
        RECT 1990.610 4.000 2008.630 4.280 ;
        RECT 2009.470 4.000 2027.950 4.280 ;
        RECT 2028.790 4.000 2046.810 4.280 ;
        RECT 2047.650 4.000 2066.130 4.280 ;
        RECT 2066.970 4.000 2084.990 4.280 ;
        RECT 2085.830 4.000 2103.850 4.280 ;
        RECT 2104.690 4.000 2123.170 4.280 ;
        RECT 2124.010 4.000 2142.030 4.280 ;
        RECT 2142.870 4.000 2161.350 4.280 ;
        RECT 2162.190 4.000 2180.210 4.280 ;
        RECT 2181.050 4.000 2199.070 4.280 ;
        RECT 2199.910 4.000 2218.390 4.280 ;
        RECT 2219.230 4.000 2237.250 4.280 ;
        RECT 2238.090 4.000 2256.570 4.280 ;
        RECT 2257.410 4.000 2275.430 4.280 ;
        RECT 2276.270 4.000 2294.290 4.280 ;
        RECT 2295.130 4.000 2313.610 4.280 ;
        RECT 2314.450 4.000 2332.470 4.280 ;
        RECT 2333.310 4.000 2351.790 4.280 ;
        RECT 2352.630 4.000 2370.650 4.280 ;
        RECT 2371.490 4.000 2389.970 4.280 ;
        RECT 2390.810 4.000 2408.830 4.280 ;
        RECT 2409.670 4.000 2427.690 4.280 ;
        RECT 2428.530 4.000 2447.010 4.280 ;
        RECT 2447.850 4.000 2465.870 4.280 ;
        RECT 2466.710 4.000 2485.190 4.280 ;
        RECT 2486.030 4.000 2504.050 4.280 ;
        RECT 2504.890 4.000 2522.910 4.280 ;
        RECT 2523.750 4.000 2542.230 4.280 ;
        RECT 2543.070 4.000 2561.090 4.280 ;
        RECT 2561.930 4.000 2580.410 4.280 ;
        RECT 2581.250 4.000 2599.270 4.280 ;
        RECT 2600.110 4.000 2618.130 4.280 ;
        RECT 2618.970 4.000 2637.450 4.280 ;
        RECT 2638.290 4.000 2656.310 4.280 ;
        RECT 2657.150 4.000 2675.630 4.280 ;
        RECT 2676.470 4.000 2694.490 4.280 ;
        RECT 2695.330 4.000 2713.350 4.280 ;
        RECT 2714.190 4.000 2732.670 4.280 ;
        RECT 2733.510 4.000 2751.530 4.280 ;
        RECT 2752.370 4.000 2770.850 4.280 ;
        RECT 2771.690 4.000 2789.710 4.280 ;
        RECT 2790.550 4.000 2791.180 4.280 ;
      LAYER met3 ;
        RECT 12.945 9.015 2790.295 688.665 ;
      LAYER met4 ;
        RECT 96.895 10.240 97.440 673.025 ;
        RECT 99.840 10.240 174.240 673.025 ;
        RECT 176.640 10.240 251.040 673.025 ;
        RECT 253.440 10.240 327.840 673.025 ;
        RECT 330.240 10.240 404.640 673.025 ;
        RECT 407.040 10.240 481.440 673.025 ;
        RECT 483.840 10.240 558.240 673.025 ;
        RECT 560.640 10.240 635.040 673.025 ;
        RECT 637.440 10.240 711.840 673.025 ;
        RECT 714.240 10.240 788.640 673.025 ;
        RECT 791.040 10.240 865.440 673.025 ;
        RECT 867.840 10.240 942.240 673.025 ;
        RECT 944.640 10.240 1019.040 673.025 ;
        RECT 1021.440 10.240 1095.840 673.025 ;
        RECT 1098.240 10.240 1172.640 673.025 ;
        RECT 1175.040 10.240 1249.440 673.025 ;
        RECT 1251.840 10.240 1326.240 673.025 ;
        RECT 1328.640 10.240 1403.040 673.025 ;
        RECT 1405.440 10.240 1479.840 673.025 ;
        RECT 1482.240 10.240 1556.640 673.025 ;
        RECT 1559.040 10.240 1633.440 673.025 ;
        RECT 1635.840 10.240 1710.240 673.025 ;
        RECT 1712.640 10.240 1787.040 673.025 ;
        RECT 1789.440 10.240 1863.840 673.025 ;
        RECT 1866.240 10.240 1940.640 673.025 ;
        RECT 1943.040 10.240 2017.440 673.025 ;
        RECT 2019.840 10.240 2094.240 673.025 ;
        RECT 2096.640 10.240 2171.040 673.025 ;
        RECT 2173.440 10.240 2247.840 673.025 ;
        RECT 2250.240 10.240 2324.640 673.025 ;
        RECT 2327.040 10.240 2401.440 673.025 ;
        RECT 2403.840 10.240 2478.240 673.025 ;
        RECT 2480.640 10.240 2555.040 673.025 ;
        RECT 2557.440 10.240 2631.840 673.025 ;
        RECT 2634.240 10.240 2708.640 673.025 ;
        RECT 2711.040 10.240 2719.225 673.025 ;
        RECT 96.895 9.015 2719.225 10.240 ;
  END
END RAM_512x64
END LIBRARY

