magic
tech sky130A
magscale 1 2
timestamp 1611815328
<< obsli1 >>
rect 1104 2159 148856 147441
<< obsm1 >>
rect 290 1300 149578 149184
<< metal2 >>
rect 386 149200 442 150000
rect 1214 149200 1270 150000
rect 2042 149200 2098 150000
rect 2962 149200 3018 150000
rect 3790 149200 3846 150000
rect 4710 149200 4766 150000
rect 5538 149200 5594 150000
rect 6366 149200 6422 150000
rect 7286 149200 7342 150000
rect 8114 149200 8170 150000
rect 9034 149200 9090 150000
rect 9862 149200 9918 150000
rect 10782 149200 10838 150000
rect 11610 149200 11666 150000
rect 12438 149200 12494 150000
rect 13358 149200 13414 150000
rect 14186 149200 14242 150000
rect 15106 149200 15162 150000
rect 15934 149200 15990 150000
rect 16854 149200 16910 150000
rect 17682 149200 17738 150000
rect 18510 149200 18566 150000
rect 19430 149200 19486 150000
rect 20258 149200 20314 150000
rect 21178 149200 21234 150000
rect 22006 149200 22062 150000
rect 22834 149200 22890 150000
rect 23754 149200 23810 150000
rect 24582 149200 24638 150000
rect 25502 149200 25558 150000
rect 26330 149200 26386 150000
rect 27250 149200 27306 150000
rect 28078 149200 28134 150000
rect 28906 149200 28962 150000
rect 29826 149200 29882 150000
rect 30654 149200 30710 150000
rect 31574 149200 31630 150000
rect 32402 149200 32458 150000
rect 33322 149200 33378 150000
rect 34150 149200 34206 150000
rect 34978 149200 35034 150000
rect 35898 149200 35954 150000
rect 36726 149200 36782 150000
rect 37646 149200 37702 150000
rect 38474 149200 38530 150000
rect 39302 149200 39358 150000
rect 40222 149200 40278 150000
rect 41050 149200 41106 150000
rect 41970 149200 42026 150000
rect 42798 149200 42854 150000
rect 43718 149200 43774 150000
rect 44546 149200 44602 150000
rect 45374 149200 45430 150000
rect 46294 149200 46350 150000
rect 47122 149200 47178 150000
rect 48042 149200 48098 150000
rect 48870 149200 48926 150000
rect 49790 149200 49846 150000
rect 50618 149200 50674 150000
rect 51446 149200 51502 150000
rect 52366 149200 52422 150000
rect 53194 149200 53250 150000
rect 54114 149200 54170 150000
rect 54942 149200 54998 150000
rect 55862 149200 55918 150000
rect 56690 149200 56746 150000
rect 57518 149200 57574 150000
rect 58438 149200 58494 150000
rect 59266 149200 59322 150000
rect 60186 149200 60242 150000
rect 61014 149200 61070 150000
rect 61842 149200 61898 150000
rect 62762 149200 62818 150000
rect 63590 149200 63646 150000
rect 64510 149200 64566 150000
rect 65338 149200 65394 150000
rect 66258 149200 66314 150000
rect 67086 149200 67142 150000
rect 67914 149200 67970 150000
rect 68834 149200 68890 150000
rect 69662 149200 69718 150000
rect 70582 149200 70638 150000
rect 71410 149200 71466 150000
rect 72330 149200 72386 150000
rect 73158 149200 73214 150000
rect 73986 149200 74042 150000
rect 74906 149200 74962 150000
rect 75734 149200 75790 150000
rect 76654 149200 76710 150000
rect 77482 149200 77538 150000
rect 78310 149200 78366 150000
rect 79230 149200 79286 150000
rect 80058 149200 80114 150000
rect 80978 149200 81034 150000
rect 81806 149200 81862 150000
rect 82726 149200 82782 150000
rect 83554 149200 83610 150000
rect 84382 149200 84438 150000
rect 85302 149200 85358 150000
rect 86130 149200 86186 150000
rect 87050 149200 87106 150000
rect 87878 149200 87934 150000
rect 88798 149200 88854 150000
rect 89626 149200 89682 150000
rect 90454 149200 90510 150000
rect 91374 149200 91430 150000
rect 92202 149200 92258 150000
rect 93122 149200 93178 150000
rect 93950 149200 94006 150000
rect 94778 149200 94834 150000
rect 95698 149200 95754 150000
rect 96526 149200 96582 150000
rect 97446 149200 97502 150000
rect 98274 149200 98330 150000
rect 99194 149200 99250 150000
rect 100022 149200 100078 150000
rect 100850 149200 100906 150000
rect 101770 149200 101826 150000
rect 102598 149200 102654 150000
rect 103518 149200 103574 150000
rect 104346 149200 104402 150000
rect 105266 149200 105322 150000
rect 106094 149200 106150 150000
rect 106922 149200 106978 150000
rect 107842 149200 107898 150000
rect 108670 149200 108726 150000
rect 109590 149200 109646 150000
rect 110418 149200 110474 150000
rect 111338 149200 111394 150000
rect 112166 149200 112222 150000
rect 112994 149200 113050 150000
rect 113914 149200 113970 150000
rect 114742 149200 114798 150000
rect 115662 149200 115718 150000
rect 116490 149200 116546 150000
rect 117318 149200 117374 150000
rect 118238 149200 118294 150000
rect 119066 149200 119122 150000
rect 119986 149200 120042 150000
rect 120814 149200 120870 150000
rect 121734 149200 121790 150000
rect 122562 149200 122618 150000
rect 123390 149200 123446 150000
rect 124310 149200 124366 150000
rect 125138 149200 125194 150000
rect 126058 149200 126114 150000
rect 126886 149200 126942 150000
rect 127806 149200 127862 150000
rect 128634 149200 128690 150000
rect 129462 149200 129518 150000
rect 130382 149200 130438 150000
rect 131210 149200 131266 150000
rect 132130 149200 132186 150000
rect 132958 149200 133014 150000
rect 133786 149200 133842 150000
rect 134706 149200 134762 150000
rect 135534 149200 135590 150000
rect 136454 149200 136510 150000
rect 137282 149200 137338 150000
rect 138202 149200 138258 150000
rect 139030 149200 139086 150000
rect 139858 149200 139914 150000
rect 140778 149200 140834 150000
rect 141606 149200 141662 150000
rect 142526 149200 142582 150000
rect 143354 149200 143410 150000
rect 144274 149200 144330 150000
rect 145102 149200 145158 150000
rect 145930 149200 145986 150000
rect 146850 149200 146906 150000
rect 147678 149200 147734 150000
rect 148598 149200 148654 150000
rect 149426 149200 149482 150000
rect 294 0 350 800
rect 938 0 994 800
rect 1674 0 1730 800
rect 2410 0 2466 800
rect 3054 0 3110 800
rect 3790 0 3846 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 8022 0 8078 800
rect 8758 0 8814 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10874 0 10930 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12990 0 13046 800
rect 13726 0 13782 800
rect 14370 0 14426 800
rect 15106 0 15162 800
rect 15842 0 15898 800
rect 16486 0 16542 800
rect 17222 0 17278 800
rect 17958 0 18014 800
rect 18602 0 18658 800
rect 19338 0 19394 800
rect 20074 0 20130 800
rect 20718 0 20774 800
rect 21454 0 21510 800
rect 22190 0 22246 800
rect 22926 0 22982 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 25042 0 25098 800
rect 25686 0 25742 800
rect 26422 0 26478 800
rect 27158 0 27214 800
rect 27802 0 27858 800
rect 28538 0 28594 800
rect 29274 0 29330 800
rect 29918 0 29974 800
rect 30654 0 30710 800
rect 31390 0 31446 800
rect 32034 0 32090 800
rect 32770 0 32826 800
rect 33506 0 33562 800
rect 34242 0 34298 800
rect 34886 0 34942 800
rect 35622 0 35678 800
rect 36358 0 36414 800
rect 37002 0 37058 800
rect 37738 0 37794 800
rect 38474 0 38530 800
rect 39118 0 39174 800
rect 39854 0 39910 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41970 0 42026 800
rect 42706 0 42762 800
rect 43442 0 43498 800
rect 44086 0 44142 800
rect 44822 0 44878 800
rect 45558 0 45614 800
rect 46202 0 46258 800
rect 46938 0 46994 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 49054 0 49110 800
rect 49790 0 49846 800
rect 50434 0 50490 800
rect 51170 0 51226 800
rect 51906 0 51962 800
rect 52550 0 52606 800
rect 53286 0 53342 800
rect 54022 0 54078 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56138 0 56194 800
rect 56874 0 56930 800
rect 57518 0 57574 800
rect 58254 0 58310 800
rect 58990 0 59046 800
rect 59634 0 59690 800
rect 60370 0 60426 800
rect 61106 0 61162 800
rect 61750 0 61806 800
rect 62486 0 62542 800
rect 63222 0 63278 800
rect 63866 0 63922 800
rect 64602 0 64658 800
rect 65338 0 65394 800
rect 66074 0 66130 800
rect 66718 0 66774 800
rect 67454 0 67510 800
rect 68190 0 68246 800
rect 68834 0 68890 800
rect 69570 0 69626 800
rect 70306 0 70362 800
rect 70950 0 71006 800
rect 71686 0 71742 800
rect 72422 0 72478 800
rect 73066 0 73122 800
rect 73802 0 73858 800
rect 74538 0 74594 800
rect 75274 0 75330 800
rect 75918 0 75974 800
rect 76654 0 76710 800
rect 77390 0 77446 800
rect 78034 0 78090 800
rect 78770 0 78826 800
rect 79506 0 79562 800
rect 80150 0 80206 800
rect 80886 0 80942 800
rect 81622 0 81678 800
rect 82266 0 82322 800
rect 83002 0 83058 800
rect 83738 0 83794 800
rect 84382 0 84438 800
rect 85118 0 85174 800
rect 85854 0 85910 800
rect 86590 0 86646 800
rect 87234 0 87290 800
rect 87970 0 88026 800
rect 88706 0 88762 800
rect 89350 0 89406 800
rect 90086 0 90142 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92202 0 92258 800
rect 92938 0 92994 800
rect 93582 0 93638 800
rect 94318 0 94374 800
rect 95054 0 95110 800
rect 95698 0 95754 800
rect 96434 0 96490 800
rect 97170 0 97226 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99286 0 99342 800
rect 100022 0 100078 800
rect 100666 0 100722 800
rect 101402 0 101458 800
rect 102138 0 102194 800
rect 102782 0 102838 800
rect 103518 0 103574 800
rect 104254 0 104310 800
rect 104898 0 104954 800
rect 105634 0 105690 800
rect 106370 0 106426 800
rect 107014 0 107070 800
rect 107750 0 107806 800
rect 108486 0 108542 800
rect 109222 0 109278 800
rect 109866 0 109922 800
rect 110602 0 110658 800
rect 111338 0 111394 800
rect 111982 0 112038 800
rect 112718 0 112774 800
rect 113454 0 113510 800
rect 114098 0 114154 800
rect 114834 0 114890 800
rect 115570 0 115626 800
rect 116214 0 116270 800
rect 116950 0 117006 800
rect 117686 0 117742 800
rect 118422 0 118478 800
rect 119066 0 119122 800
rect 119802 0 119858 800
rect 120538 0 120594 800
rect 121182 0 121238 800
rect 121918 0 121974 800
rect 122654 0 122710 800
rect 123298 0 123354 800
rect 124034 0 124090 800
rect 124770 0 124826 800
rect 125414 0 125470 800
rect 126150 0 126206 800
rect 126886 0 126942 800
rect 127530 0 127586 800
rect 128266 0 128322 800
rect 129002 0 129058 800
rect 129738 0 129794 800
rect 130382 0 130438 800
rect 131118 0 131174 800
rect 131854 0 131910 800
rect 132498 0 132554 800
rect 133234 0 133290 800
rect 133970 0 134026 800
rect 134614 0 134670 800
rect 135350 0 135406 800
rect 136086 0 136142 800
rect 136730 0 136786 800
rect 137466 0 137522 800
rect 138202 0 138258 800
rect 138846 0 138902 800
rect 139582 0 139638 800
rect 140318 0 140374 800
rect 141054 0 141110 800
rect 141698 0 141754 800
rect 142434 0 142490 800
rect 143170 0 143226 800
rect 143814 0 143870 800
rect 144550 0 144606 800
rect 145286 0 145342 800
rect 145930 0 145986 800
rect 146666 0 146722 800
rect 147402 0 147458 800
rect 148046 0 148102 800
rect 148782 0 148838 800
rect 149518 0 149574 800
<< obsm2 >>
rect 296 149144 330 149569
rect 498 149144 1158 149569
rect 1326 149144 1986 149569
rect 2154 149144 2906 149569
rect 3074 149144 3734 149569
rect 3902 149144 4654 149569
rect 4822 149144 5482 149569
rect 5650 149144 6310 149569
rect 6478 149144 7230 149569
rect 7398 149144 8058 149569
rect 8226 149144 8978 149569
rect 9146 149144 9806 149569
rect 9974 149144 10726 149569
rect 10894 149144 11554 149569
rect 11722 149144 12382 149569
rect 12550 149144 13302 149569
rect 13470 149144 14130 149569
rect 14298 149144 15050 149569
rect 15218 149144 15878 149569
rect 16046 149144 16798 149569
rect 16966 149144 17626 149569
rect 17794 149144 18454 149569
rect 18622 149144 19374 149569
rect 19542 149144 20202 149569
rect 20370 149144 21122 149569
rect 21290 149144 21950 149569
rect 22118 149144 22778 149569
rect 22946 149144 23698 149569
rect 23866 149144 24526 149569
rect 24694 149144 25446 149569
rect 25614 149144 26274 149569
rect 26442 149144 27194 149569
rect 27362 149144 28022 149569
rect 28190 149144 28850 149569
rect 29018 149144 29770 149569
rect 29938 149144 30598 149569
rect 30766 149144 31518 149569
rect 31686 149144 32346 149569
rect 32514 149144 33266 149569
rect 33434 149144 34094 149569
rect 34262 149144 34922 149569
rect 35090 149144 35842 149569
rect 36010 149144 36670 149569
rect 36838 149144 37590 149569
rect 37758 149144 38418 149569
rect 38586 149144 39246 149569
rect 39414 149144 40166 149569
rect 40334 149144 40994 149569
rect 41162 149144 41914 149569
rect 42082 149144 42742 149569
rect 42910 149144 43662 149569
rect 43830 149144 44490 149569
rect 44658 149144 45318 149569
rect 45486 149144 46238 149569
rect 46406 149144 47066 149569
rect 47234 149144 47986 149569
rect 48154 149144 48814 149569
rect 48982 149144 49734 149569
rect 49902 149144 50562 149569
rect 50730 149144 51390 149569
rect 51558 149144 52310 149569
rect 52478 149144 53138 149569
rect 53306 149144 54058 149569
rect 54226 149144 54886 149569
rect 55054 149144 55806 149569
rect 55974 149144 56634 149569
rect 56802 149144 57462 149569
rect 57630 149144 58382 149569
rect 58550 149144 59210 149569
rect 59378 149144 60130 149569
rect 60298 149144 60958 149569
rect 61126 149144 61786 149569
rect 61954 149144 62706 149569
rect 62874 149144 63534 149569
rect 63702 149144 64454 149569
rect 64622 149144 65282 149569
rect 65450 149144 66202 149569
rect 66370 149144 67030 149569
rect 67198 149144 67858 149569
rect 68026 149144 68778 149569
rect 68946 149144 69606 149569
rect 69774 149144 70526 149569
rect 70694 149144 71354 149569
rect 71522 149144 72274 149569
rect 72442 149144 73102 149569
rect 73270 149144 73930 149569
rect 74098 149144 74850 149569
rect 75018 149144 75678 149569
rect 75846 149144 76598 149569
rect 76766 149144 77426 149569
rect 77594 149144 78254 149569
rect 78422 149144 79174 149569
rect 79342 149144 80002 149569
rect 80170 149144 80922 149569
rect 81090 149144 81750 149569
rect 81918 149144 82670 149569
rect 82838 149144 83498 149569
rect 83666 149144 84326 149569
rect 84494 149144 85246 149569
rect 85414 149144 86074 149569
rect 86242 149144 86994 149569
rect 87162 149144 87822 149569
rect 87990 149144 88742 149569
rect 88910 149144 89570 149569
rect 89738 149144 90398 149569
rect 90566 149144 91318 149569
rect 91486 149144 92146 149569
rect 92314 149144 93066 149569
rect 93234 149144 93894 149569
rect 94062 149144 94722 149569
rect 94890 149144 95642 149569
rect 95810 149144 96470 149569
rect 96638 149144 97390 149569
rect 97558 149144 98218 149569
rect 98386 149144 99138 149569
rect 99306 149144 99966 149569
rect 100134 149144 100794 149569
rect 100962 149144 101714 149569
rect 101882 149144 102542 149569
rect 102710 149144 103462 149569
rect 103630 149144 104290 149569
rect 104458 149144 105210 149569
rect 105378 149144 106038 149569
rect 106206 149144 106866 149569
rect 107034 149144 107786 149569
rect 107954 149144 108614 149569
rect 108782 149144 109534 149569
rect 109702 149144 110362 149569
rect 110530 149144 111282 149569
rect 111450 149144 112110 149569
rect 112278 149144 112938 149569
rect 113106 149144 113858 149569
rect 114026 149144 114686 149569
rect 114854 149144 115606 149569
rect 115774 149144 116434 149569
rect 116602 149144 117262 149569
rect 117430 149144 118182 149569
rect 118350 149144 119010 149569
rect 119178 149144 119930 149569
rect 120098 149144 120758 149569
rect 120926 149144 121678 149569
rect 121846 149144 122506 149569
rect 122674 149144 123334 149569
rect 123502 149144 124254 149569
rect 124422 149144 125082 149569
rect 125250 149144 126002 149569
rect 126170 149144 126830 149569
rect 126998 149144 127750 149569
rect 127918 149144 128578 149569
rect 128746 149144 129406 149569
rect 129574 149144 130326 149569
rect 130494 149144 131154 149569
rect 131322 149144 132074 149569
rect 132242 149144 132902 149569
rect 133070 149144 133730 149569
rect 133898 149144 134650 149569
rect 134818 149144 135478 149569
rect 135646 149144 136398 149569
rect 136566 149144 137226 149569
rect 137394 149144 138146 149569
rect 138314 149144 138974 149569
rect 139142 149144 139802 149569
rect 139970 149144 140722 149569
rect 140890 149144 141550 149569
rect 141718 149144 142470 149569
rect 142638 149144 143298 149569
rect 143466 149144 144218 149569
rect 144386 149144 145046 149569
rect 145214 149144 145874 149569
rect 146042 149144 146794 149569
rect 146962 149144 147622 149569
rect 147790 149144 148542 149569
rect 148710 149144 149370 149569
rect 149538 149144 149572 149569
rect 296 856 149572 149144
rect 406 303 882 856
rect 1050 303 1618 856
rect 1786 303 2354 856
rect 2522 303 2998 856
rect 3166 303 3734 856
rect 3902 303 4470 856
rect 4638 303 5114 856
rect 5282 303 5850 856
rect 6018 303 6586 856
rect 6754 303 7230 856
rect 7398 303 7966 856
rect 8134 303 8702 856
rect 8870 303 9346 856
rect 9514 303 10082 856
rect 10250 303 10818 856
rect 10986 303 11554 856
rect 11722 303 12198 856
rect 12366 303 12934 856
rect 13102 303 13670 856
rect 13838 303 14314 856
rect 14482 303 15050 856
rect 15218 303 15786 856
rect 15954 303 16430 856
rect 16598 303 17166 856
rect 17334 303 17902 856
rect 18070 303 18546 856
rect 18714 303 19282 856
rect 19450 303 20018 856
rect 20186 303 20662 856
rect 20830 303 21398 856
rect 21566 303 22134 856
rect 22302 303 22870 856
rect 23038 303 23514 856
rect 23682 303 24250 856
rect 24418 303 24986 856
rect 25154 303 25630 856
rect 25798 303 26366 856
rect 26534 303 27102 856
rect 27270 303 27746 856
rect 27914 303 28482 856
rect 28650 303 29218 856
rect 29386 303 29862 856
rect 30030 303 30598 856
rect 30766 303 31334 856
rect 31502 303 31978 856
rect 32146 303 32714 856
rect 32882 303 33450 856
rect 33618 303 34186 856
rect 34354 303 34830 856
rect 34998 303 35566 856
rect 35734 303 36302 856
rect 36470 303 36946 856
rect 37114 303 37682 856
rect 37850 303 38418 856
rect 38586 303 39062 856
rect 39230 303 39798 856
rect 39966 303 40534 856
rect 40702 303 41178 856
rect 41346 303 41914 856
rect 42082 303 42650 856
rect 42818 303 43386 856
rect 43554 303 44030 856
rect 44198 303 44766 856
rect 44934 303 45502 856
rect 45670 303 46146 856
rect 46314 303 46882 856
rect 47050 303 47618 856
rect 47786 303 48262 856
rect 48430 303 48998 856
rect 49166 303 49734 856
rect 49902 303 50378 856
rect 50546 303 51114 856
rect 51282 303 51850 856
rect 52018 303 52494 856
rect 52662 303 53230 856
rect 53398 303 53966 856
rect 54134 303 54702 856
rect 54870 303 55346 856
rect 55514 303 56082 856
rect 56250 303 56818 856
rect 56986 303 57462 856
rect 57630 303 58198 856
rect 58366 303 58934 856
rect 59102 303 59578 856
rect 59746 303 60314 856
rect 60482 303 61050 856
rect 61218 303 61694 856
rect 61862 303 62430 856
rect 62598 303 63166 856
rect 63334 303 63810 856
rect 63978 303 64546 856
rect 64714 303 65282 856
rect 65450 303 66018 856
rect 66186 303 66662 856
rect 66830 303 67398 856
rect 67566 303 68134 856
rect 68302 303 68778 856
rect 68946 303 69514 856
rect 69682 303 70250 856
rect 70418 303 70894 856
rect 71062 303 71630 856
rect 71798 303 72366 856
rect 72534 303 73010 856
rect 73178 303 73746 856
rect 73914 303 74482 856
rect 74650 303 75218 856
rect 75386 303 75862 856
rect 76030 303 76598 856
rect 76766 303 77334 856
rect 77502 303 77978 856
rect 78146 303 78714 856
rect 78882 303 79450 856
rect 79618 303 80094 856
rect 80262 303 80830 856
rect 80998 303 81566 856
rect 81734 303 82210 856
rect 82378 303 82946 856
rect 83114 303 83682 856
rect 83850 303 84326 856
rect 84494 303 85062 856
rect 85230 303 85798 856
rect 85966 303 86534 856
rect 86702 303 87178 856
rect 87346 303 87914 856
rect 88082 303 88650 856
rect 88818 303 89294 856
rect 89462 303 90030 856
rect 90198 303 90766 856
rect 90934 303 91410 856
rect 91578 303 92146 856
rect 92314 303 92882 856
rect 93050 303 93526 856
rect 93694 303 94262 856
rect 94430 303 94998 856
rect 95166 303 95642 856
rect 95810 303 96378 856
rect 96546 303 97114 856
rect 97282 303 97850 856
rect 98018 303 98494 856
rect 98662 303 99230 856
rect 99398 303 99966 856
rect 100134 303 100610 856
rect 100778 303 101346 856
rect 101514 303 102082 856
rect 102250 303 102726 856
rect 102894 303 103462 856
rect 103630 303 104198 856
rect 104366 303 104842 856
rect 105010 303 105578 856
rect 105746 303 106314 856
rect 106482 303 106958 856
rect 107126 303 107694 856
rect 107862 303 108430 856
rect 108598 303 109166 856
rect 109334 303 109810 856
rect 109978 303 110546 856
rect 110714 303 111282 856
rect 111450 303 111926 856
rect 112094 303 112662 856
rect 112830 303 113398 856
rect 113566 303 114042 856
rect 114210 303 114778 856
rect 114946 303 115514 856
rect 115682 303 116158 856
rect 116326 303 116894 856
rect 117062 303 117630 856
rect 117798 303 118366 856
rect 118534 303 119010 856
rect 119178 303 119746 856
rect 119914 303 120482 856
rect 120650 303 121126 856
rect 121294 303 121862 856
rect 122030 303 122598 856
rect 122766 303 123242 856
rect 123410 303 123978 856
rect 124146 303 124714 856
rect 124882 303 125358 856
rect 125526 303 126094 856
rect 126262 303 126830 856
rect 126998 303 127474 856
rect 127642 303 128210 856
rect 128378 303 128946 856
rect 129114 303 129682 856
rect 129850 303 130326 856
rect 130494 303 131062 856
rect 131230 303 131798 856
rect 131966 303 132442 856
rect 132610 303 133178 856
rect 133346 303 133914 856
rect 134082 303 134558 856
rect 134726 303 135294 856
rect 135462 303 136030 856
rect 136198 303 136674 856
rect 136842 303 137410 856
rect 137578 303 138146 856
rect 138314 303 138790 856
rect 138958 303 139526 856
rect 139694 303 140262 856
rect 140430 303 140998 856
rect 141166 303 141642 856
rect 141810 303 142378 856
rect 142546 303 143114 856
rect 143282 303 143758 856
rect 143926 303 144494 856
rect 144662 303 145230 856
rect 145398 303 145874 856
rect 146042 303 146610 856
rect 146778 303 147346 856
rect 147514 303 147990 856
rect 148158 303 148726 856
rect 148894 303 149462 856
<< metal3 >>
rect 0 149472 800 149592
rect 0 148792 800 148912
rect 0 147976 800 148096
rect 0 147296 800 147416
rect 0 146480 800 146600
rect 0 145800 800 145920
rect 0 144984 800 145104
rect 0 144304 800 144424
rect 0 143488 800 143608
rect 0 142808 800 142928
rect 0 141992 800 142112
rect 0 141312 800 141432
rect 0 140496 800 140616
rect 0 139816 800 139936
rect 0 139000 800 139120
rect 0 138320 800 138440
rect 0 137504 800 137624
rect 0 136824 800 136944
rect 0 136008 800 136128
rect 0 135328 800 135448
rect 0 134512 800 134632
rect 0 133832 800 133952
rect 0 133016 800 133136
rect 0 132336 800 132456
rect 0 131520 800 131640
rect 0 130840 800 130960
rect 0 130024 800 130144
rect 0 129344 800 129464
rect 0 128528 800 128648
rect 0 127848 800 127968
rect 0 127032 800 127152
rect 0 126352 800 126472
rect 0 125536 800 125656
rect 0 124856 800 124976
rect 0 124040 800 124160
rect 0 123360 800 123480
rect 0 122544 800 122664
rect 0 121864 800 121984
rect 0 121048 800 121168
rect 0 120368 800 120488
rect 0 119688 800 119808
rect 0 118872 800 118992
rect 0 118192 800 118312
rect 0 117376 800 117496
rect 0 116696 800 116816
rect 0 115880 800 116000
rect 0 115200 800 115320
rect 0 114384 800 114504
rect 0 113704 800 113824
rect 0 112888 800 113008
rect 0 112208 800 112328
rect 0 111392 800 111512
rect 0 110712 800 110832
rect 0 109896 800 110016
rect 0 109216 800 109336
rect 0 108400 800 108520
rect 0 107720 800 107840
rect 0 106904 800 107024
rect 0 106224 800 106344
rect 0 105408 800 105528
rect 0 104728 800 104848
rect 0 103912 800 104032
rect 0 103232 800 103352
rect 0 102416 800 102536
rect 0 101736 800 101856
rect 0 100920 800 101040
rect 0 100240 800 100360
rect 0 99424 800 99544
rect 0 98744 800 98864
rect 0 97928 800 98048
rect 0 97248 800 97368
rect 0 96432 800 96552
rect 0 95752 800 95872
rect 0 94936 800 95056
rect 0 94256 800 94376
rect 0 93440 800 93560
rect 0 92760 800 92880
rect 0 91944 800 92064
rect 0 91264 800 91384
rect 0 90448 800 90568
rect 0 89768 800 89888
rect 0 89088 800 89208
rect 0 88272 800 88392
rect 0 87592 800 87712
rect 0 86776 800 86896
rect 0 86096 800 86216
rect 0 85280 800 85400
rect 0 84600 800 84720
rect 0 83784 800 83904
rect 0 83104 800 83224
rect 0 82288 800 82408
rect 0 81608 800 81728
rect 0 80792 800 80912
rect 0 80112 800 80232
rect 0 79296 800 79416
rect 0 78616 800 78736
rect 0 77800 800 77920
rect 0 77120 800 77240
rect 0 76304 800 76424
rect 0 75624 800 75744
rect 0 74808 800 74928
rect 0 74128 800 74248
rect 0 73312 800 73432
rect 0 72632 800 72752
rect 0 71816 800 71936
rect 0 71136 800 71256
rect 0 70320 800 70440
rect 0 69640 800 69760
rect 0 68824 800 68944
rect 0 68144 800 68264
rect 0 67328 800 67448
rect 0 66648 800 66768
rect 0 65832 800 65952
rect 0 65152 800 65272
rect 0 64336 800 64456
rect 0 63656 800 63776
rect 0 62840 800 62960
rect 0 62160 800 62280
rect 0 61344 800 61464
rect 0 60664 800 60784
rect 0 59984 800 60104
rect 0 59168 800 59288
rect 0 58488 800 58608
rect 0 57672 800 57792
rect 0 56992 800 57112
rect 0 56176 800 56296
rect 0 55496 800 55616
rect 0 54680 800 54800
rect 0 54000 800 54120
rect 0 53184 800 53304
rect 0 52504 800 52624
rect 0 51688 800 51808
rect 0 51008 800 51128
rect 0 50192 800 50312
rect 0 49512 800 49632
rect 0 48696 800 48816
rect 0 48016 800 48136
rect 0 47200 800 47320
rect 0 46520 800 46640
rect 0 45704 800 45824
rect 0 45024 800 45144
rect 0 44208 800 44328
rect 0 43528 800 43648
rect 0 42712 800 42832
rect 0 42032 800 42152
rect 0 41216 800 41336
rect 0 40536 800 40656
rect 0 39720 800 39840
rect 0 39040 800 39160
rect 0 38224 800 38344
rect 0 37544 800 37664
rect 0 36728 800 36848
rect 0 36048 800 36168
rect 0 35232 800 35352
rect 0 34552 800 34672
rect 0 33736 800 33856
rect 0 33056 800 33176
rect 0 32240 800 32360
rect 0 31560 800 31680
rect 0 30744 800 30864
rect 0 30064 800 30184
rect 0 29384 800 29504
rect 0 28568 800 28688
rect 0 27888 800 28008
rect 0 27072 800 27192
rect 0 26392 800 26512
rect 0 25576 800 25696
rect 0 24896 800 25016
rect 0 24080 800 24200
rect 0 23400 800 23520
rect 0 22584 800 22704
rect 0 21904 800 22024
rect 0 21088 800 21208
rect 0 20408 800 20528
rect 0 19592 800 19712
rect 0 18912 800 19032
rect 0 18096 800 18216
rect 0 17416 800 17536
rect 0 16600 800 16720
rect 0 15920 800 16040
rect 0 15104 800 15224
rect 0 14424 800 14544
rect 0 13608 800 13728
rect 0 12928 800 13048
rect 0 12112 800 12232
rect 0 11432 800 11552
rect 0 10616 800 10736
rect 0 9936 800 10056
rect 0 9120 800 9240
rect 0 8440 800 8560
rect 0 7624 800 7744
rect 0 6944 800 7064
rect 0 6128 800 6248
rect 0 5448 800 5568
rect 0 4632 800 4752
rect 0 3952 800 4072
rect 0 3136 800 3256
rect 0 2456 800 2576
rect 0 1640 800 1760
rect 0 960 800 1080
rect 0 280 800 400
<< obsm3 >>
rect 880 149392 148383 149565
rect 238 148992 148383 149392
rect 880 148712 148383 148992
rect 238 148176 148383 148712
rect 880 147896 148383 148176
rect 238 147496 148383 147896
rect 880 147216 148383 147496
rect 238 146680 148383 147216
rect 880 146400 148383 146680
rect 238 146000 148383 146400
rect 880 145720 148383 146000
rect 238 145184 148383 145720
rect 880 144904 148383 145184
rect 238 144504 148383 144904
rect 880 144224 148383 144504
rect 238 143688 148383 144224
rect 880 143408 148383 143688
rect 238 143008 148383 143408
rect 880 142728 148383 143008
rect 238 142192 148383 142728
rect 880 141912 148383 142192
rect 238 141512 148383 141912
rect 880 141232 148383 141512
rect 238 140696 148383 141232
rect 880 140416 148383 140696
rect 238 140016 148383 140416
rect 880 139736 148383 140016
rect 238 139200 148383 139736
rect 880 138920 148383 139200
rect 238 138520 148383 138920
rect 880 138240 148383 138520
rect 238 137704 148383 138240
rect 880 137424 148383 137704
rect 238 137024 148383 137424
rect 880 136744 148383 137024
rect 238 136208 148383 136744
rect 880 135928 148383 136208
rect 238 135528 148383 135928
rect 880 135248 148383 135528
rect 238 134712 148383 135248
rect 880 134432 148383 134712
rect 238 134032 148383 134432
rect 880 133752 148383 134032
rect 238 133216 148383 133752
rect 880 132936 148383 133216
rect 238 132536 148383 132936
rect 880 132256 148383 132536
rect 238 131720 148383 132256
rect 880 131440 148383 131720
rect 238 131040 148383 131440
rect 880 130760 148383 131040
rect 238 130224 148383 130760
rect 880 129944 148383 130224
rect 238 129544 148383 129944
rect 880 129264 148383 129544
rect 238 128728 148383 129264
rect 880 128448 148383 128728
rect 238 128048 148383 128448
rect 880 127768 148383 128048
rect 238 127232 148383 127768
rect 880 126952 148383 127232
rect 238 126552 148383 126952
rect 880 126272 148383 126552
rect 238 125736 148383 126272
rect 880 125456 148383 125736
rect 238 125056 148383 125456
rect 880 124776 148383 125056
rect 238 124240 148383 124776
rect 880 123960 148383 124240
rect 238 123560 148383 123960
rect 880 123280 148383 123560
rect 238 122744 148383 123280
rect 880 122464 148383 122744
rect 238 122064 148383 122464
rect 880 121784 148383 122064
rect 238 121248 148383 121784
rect 880 120968 148383 121248
rect 238 120568 148383 120968
rect 880 120288 148383 120568
rect 238 119888 148383 120288
rect 880 119608 148383 119888
rect 238 119072 148383 119608
rect 880 118792 148383 119072
rect 238 118392 148383 118792
rect 880 118112 148383 118392
rect 238 117576 148383 118112
rect 880 117296 148383 117576
rect 238 116896 148383 117296
rect 880 116616 148383 116896
rect 238 116080 148383 116616
rect 880 115800 148383 116080
rect 238 115400 148383 115800
rect 880 115120 148383 115400
rect 238 114584 148383 115120
rect 880 114304 148383 114584
rect 238 113904 148383 114304
rect 880 113624 148383 113904
rect 238 113088 148383 113624
rect 880 112808 148383 113088
rect 238 112408 148383 112808
rect 880 112128 148383 112408
rect 238 111592 148383 112128
rect 880 111312 148383 111592
rect 238 110912 148383 111312
rect 880 110632 148383 110912
rect 238 110096 148383 110632
rect 880 109816 148383 110096
rect 238 109416 148383 109816
rect 880 109136 148383 109416
rect 238 108600 148383 109136
rect 880 108320 148383 108600
rect 238 107920 148383 108320
rect 880 107640 148383 107920
rect 238 107104 148383 107640
rect 880 106824 148383 107104
rect 238 106424 148383 106824
rect 880 106144 148383 106424
rect 238 105608 148383 106144
rect 880 105328 148383 105608
rect 238 104928 148383 105328
rect 880 104648 148383 104928
rect 238 104112 148383 104648
rect 880 103832 148383 104112
rect 238 103432 148383 103832
rect 880 103152 148383 103432
rect 238 102616 148383 103152
rect 880 102336 148383 102616
rect 238 101936 148383 102336
rect 880 101656 148383 101936
rect 238 101120 148383 101656
rect 880 100840 148383 101120
rect 238 100440 148383 100840
rect 880 100160 148383 100440
rect 238 99624 148383 100160
rect 880 99344 148383 99624
rect 238 98944 148383 99344
rect 880 98664 148383 98944
rect 238 98128 148383 98664
rect 880 97848 148383 98128
rect 238 97448 148383 97848
rect 880 97168 148383 97448
rect 238 96632 148383 97168
rect 880 96352 148383 96632
rect 238 95952 148383 96352
rect 880 95672 148383 95952
rect 238 95136 148383 95672
rect 880 94856 148383 95136
rect 238 94456 148383 94856
rect 880 94176 148383 94456
rect 238 93640 148383 94176
rect 880 93360 148383 93640
rect 238 92960 148383 93360
rect 880 92680 148383 92960
rect 238 92144 148383 92680
rect 880 91864 148383 92144
rect 238 91464 148383 91864
rect 880 91184 148383 91464
rect 238 90648 148383 91184
rect 880 90368 148383 90648
rect 238 89968 148383 90368
rect 880 89688 148383 89968
rect 238 89288 148383 89688
rect 880 89008 148383 89288
rect 238 88472 148383 89008
rect 880 88192 148383 88472
rect 238 87792 148383 88192
rect 880 87512 148383 87792
rect 238 86976 148383 87512
rect 880 86696 148383 86976
rect 238 86296 148383 86696
rect 880 86016 148383 86296
rect 238 85480 148383 86016
rect 880 85200 148383 85480
rect 238 84800 148383 85200
rect 880 84520 148383 84800
rect 238 83984 148383 84520
rect 880 83704 148383 83984
rect 238 83304 148383 83704
rect 880 83024 148383 83304
rect 238 82488 148383 83024
rect 880 82208 148383 82488
rect 238 81808 148383 82208
rect 880 81528 148383 81808
rect 238 80992 148383 81528
rect 880 80712 148383 80992
rect 238 80312 148383 80712
rect 880 80032 148383 80312
rect 238 79496 148383 80032
rect 880 79216 148383 79496
rect 238 78816 148383 79216
rect 880 78536 148383 78816
rect 238 78000 148383 78536
rect 880 77720 148383 78000
rect 238 77320 148383 77720
rect 880 77040 148383 77320
rect 238 76504 148383 77040
rect 880 76224 148383 76504
rect 238 75824 148383 76224
rect 880 75544 148383 75824
rect 238 75008 148383 75544
rect 880 74728 148383 75008
rect 238 74328 148383 74728
rect 880 74048 148383 74328
rect 238 73512 148383 74048
rect 880 73232 148383 73512
rect 238 72832 148383 73232
rect 880 72552 148383 72832
rect 238 72016 148383 72552
rect 880 71736 148383 72016
rect 238 71336 148383 71736
rect 880 71056 148383 71336
rect 238 70520 148383 71056
rect 880 70240 148383 70520
rect 238 69840 148383 70240
rect 880 69560 148383 69840
rect 238 69024 148383 69560
rect 880 68744 148383 69024
rect 238 68344 148383 68744
rect 880 68064 148383 68344
rect 238 67528 148383 68064
rect 880 67248 148383 67528
rect 238 66848 148383 67248
rect 880 66568 148383 66848
rect 238 66032 148383 66568
rect 880 65752 148383 66032
rect 238 65352 148383 65752
rect 880 65072 148383 65352
rect 238 64536 148383 65072
rect 880 64256 148383 64536
rect 238 63856 148383 64256
rect 880 63576 148383 63856
rect 238 63040 148383 63576
rect 880 62760 148383 63040
rect 238 62360 148383 62760
rect 880 62080 148383 62360
rect 238 61544 148383 62080
rect 880 61264 148383 61544
rect 238 60864 148383 61264
rect 880 60584 148383 60864
rect 238 60184 148383 60584
rect 880 59904 148383 60184
rect 238 59368 148383 59904
rect 880 59088 148383 59368
rect 238 58688 148383 59088
rect 880 58408 148383 58688
rect 238 57872 148383 58408
rect 880 57592 148383 57872
rect 238 57192 148383 57592
rect 880 56912 148383 57192
rect 238 56376 148383 56912
rect 880 56096 148383 56376
rect 238 55696 148383 56096
rect 880 55416 148383 55696
rect 238 54880 148383 55416
rect 880 54600 148383 54880
rect 238 54200 148383 54600
rect 880 53920 148383 54200
rect 238 53384 148383 53920
rect 880 53104 148383 53384
rect 238 52704 148383 53104
rect 880 52424 148383 52704
rect 238 51888 148383 52424
rect 880 51608 148383 51888
rect 238 51208 148383 51608
rect 880 50928 148383 51208
rect 238 50392 148383 50928
rect 880 50112 148383 50392
rect 238 49712 148383 50112
rect 880 49432 148383 49712
rect 238 48896 148383 49432
rect 880 48616 148383 48896
rect 238 48216 148383 48616
rect 880 47936 148383 48216
rect 238 47400 148383 47936
rect 880 47120 148383 47400
rect 238 46720 148383 47120
rect 880 46440 148383 46720
rect 238 45904 148383 46440
rect 880 45624 148383 45904
rect 238 45224 148383 45624
rect 880 44944 148383 45224
rect 238 44408 148383 44944
rect 880 44128 148383 44408
rect 238 43728 148383 44128
rect 880 43448 148383 43728
rect 238 42912 148383 43448
rect 880 42632 148383 42912
rect 238 42232 148383 42632
rect 880 41952 148383 42232
rect 238 41416 148383 41952
rect 880 41136 148383 41416
rect 238 40736 148383 41136
rect 880 40456 148383 40736
rect 238 39920 148383 40456
rect 880 39640 148383 39920
rect 238 39240 148383 39640
rect 880 38960 148383 39240
rect 238 38424 148383 38960
rect 880 38144 148383 38424
rect 238 37744 148383 38144
rect 880 37464 148383 37744
rect 238 36928 148383 37464
rect 880 36648 148383 36928
rect 238 36248 148383 36648
rect 880 35968 148383 36248
rect 238 35432 148383 35968
rect 880 35152 148383 35432
rect 238 34752 148383 35152
rect 880 34472 148383 34752
rect 238 33936 148383 34472
rect 880 33656 148383 33936
rect 238 33256 148383 33656
rect 880 32976 148383 33256
rect 238 32440 148383 32976
rect 880 32160 148383 32440
rect 238 31760 148383 32160
rect 880 31480 148383 31760
rect 238 30944 148383 31480
rect 880 30664 148383 30944
rect 238 30264 148383 30664
rect 880 29984 148383 30264
rect 238 29584 148383 29984
rect 880 29304 148383 29584
rect 238 28768 148383 29304
rect 880 28488 148383 28768
rect 238 28088 148383 28488
rect 880 27808 148383 28088
rect 238 27272 148383 27808
rect 880 26992 148383 27272
rect 238 26592 148383 26992
rect 880 26312 148383 26592
rect 238 25776 148383 26312
rect 880 25496 148383 25776
rect 238 25096 148383 25496
rect 880 24816 148383 25096
rect 238 24280 148383 24816
rect 880 24000 148383 24280
rect 238 23600 148383 24000
rect 880 23320 148383 23600
rect 238 22784 148383 23320
rect 880 22504 148383 22784
rect 238 22104 148383 22504
rect 880 21824 148383 22104
rect 238 21288 148383 21824
rect 880 21008 148383 21288
rect 238 20608 148383 21008
rect 880 20328 148383 20608
rect 238 19792 148383 20328
rect 880 19512 148383 19792
rect 238 19112 148383 19512
rect 880 18832 148383 19112
rect 238 18296 148383 18832
rect 880 18016 148383 18296
rect 238 17616 148383 18016
rect 880 17336 148383 17616
rect 238 16800 148383 17336
rect 880 16520 148383 16800
rect 238 16120 148383 16520
rect 880 15840 148383 16120
rect 238 15304 148383 15840
rect 880 15024 148383 15304
rect 238 14624 148383 15024
rect 880 14344 148383 14624
rect 238 13808 148383 14344
rect 880 13528 148383 13808
rect 238 13128 148383 13528
rect 880 12848 148383 13128
rect 238 12312 148383 12848
rect 880 12032 148383 12312
rect 238 11632 148383 12032
rect 880 11352 148383 11632
rect 238 10816 148383 11352
rect 880 10536 148383 10816
rect 238 10136 148383 10536
rect 880 9856 148383 10136
rect 238 9320 148383 9856
rect 880 9040 148383 9320
rect 238 8640 148383 9040
rect 880 8360 148383 8640
rect 238 7824 148383 8360
rect 880 7544 148383 7824
rect 238 7144 148383 7544
rect 880 6864 148383 7144
rect 238 6328 148383 6864
rect 880 6048 148383 6328
rect 238 5648 148383 6048
rect 880 5368 148383 5648
rect 238 4832 148383 5368
rect 880 4552 148383 4832
rect 238 4152 148383 4552
rect 880 3872 148383 4152
rect 238 3336 148383 3872
rect 880 3056 148383 3336
rect 238 2656 148383 3056
rect 880 2376 148383 2656
rect 238 1840 148383 2376
rect 880 1560 148383 1840
rect 238 1160 148383 1560
rect 880 880 148383 1160
rect 238 480 148383 880
rect 880 307 148383 480
<< metal4 >>
rect 4208 2128 4528 147472
rect 19568 2128 19888 147472
rect 34928 2128 35248 147472
rect 50288 2128 50608 147472
rect 65648 2128 65968 147472
rect 81008 2128 81328 147472
rect 96368 2128 96688 147472
rect 111728 2128 112048 147472
rect 127088 2128 127408 147472
rect 142448 2128 142768 147472
<< obsm4 >>
rect 243 147552 146589 147797
rect 243 2048 4128 147552
rect 4608 2048 19488 147552
rect 19968 2048 34848 147552
rect 35328 2048 50208 147552
rect 50688 2048 65568 147552
rect 66048 2048 80928 147552
rect 81408 2048 96288 147552
rect 96768 2048 111648 147552
rect 112128 2048 127008 147552
rect 127488 2048 142368 147552
rect 142848 2048 146589 147552
rect 243 1259 146589 2048
<< labels >>
rlabel metal3 s 0 280 800 400 6 clk
port 1 nsew signal input
rlabel metal2 s 938 0 994 800 6 d_in[0]
port 2 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 d_in[100]
port 3 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 d_in[101]
port 4 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 d_in[102]
port 5 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 d_in[103]
port 6 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 d_in[104]
port 7 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 d_in[105]
port 8 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 d_in[106]
port 9 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 d_in[107]
port 10 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 d_in[108]
port 11 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 d_in[109]
port 12 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 d_in[10]
port 13 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 d_in[110]
port 14 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 d_in[111]
port 15 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 d_in[112]
port 16 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 d_in[113]
port 17 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 d_in[114]
port 18 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 d_in[115]
port 19 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 d_in[116]
port 20 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 d_in[117]
port 21 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 d_in[118]
port 22 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 d_in[119]
port 23 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 d_in[11]
port 24 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 d_in[120]
port 25 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 d_in[121]
port 26 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 d_in[122]
port 27 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 d_in[123]
port 28 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 d_in[124]
port 29 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 d_in[125]
port 30 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 d_in[126]
port 31 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 d_in[127]
port 32 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 d_in[128]
port 33 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 d_in[129]
port 34 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 d_in[12]
port 35 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 d_in[130]
port 36 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 d_in[131]
port 37 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 d_in[132]
port 38 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 d_in[133]
port 39 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 d_in[134]
port 40 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 d_in[135]
port 41 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 d_in[136]
port 42 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 d_in[137]
port 43 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 d_in[138]
port 44 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 d_in[139]
port 45 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 d_in[13]
port 46 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 d_in[140]
port 47 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 d_in[141]
port 48 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 d_in[142]
port 49 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 d_in[14]
port 50 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 d_in[15]
port 51 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 d_in[16]
port 52 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 d_in[17]
port 53 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 d_in[18]
port 54 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 d_in[19]
port 55 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 d_in[1]
port 56 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 d_in[20]
port 57 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 d_in[21]
port 58 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 d_in[22]
port 59 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 d_in[23]
port 60 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 d_in[24]
port 61 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 d_in[25]
port 62 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 d_in[26]
port 63 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 d_in[27]
port 64 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 d_in[28]
port 65 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 d_in[29]
port 66 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 d_in[2]
port 67 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 d_in[30]
port 68 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 d_in[31]
port 69 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 d_in[32]
port 70 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 d_in[33]
port 71 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 d_in[34]
port 72 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 d_in[35]
port 73 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 d_in[36]
port 74 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 d_in[37]
port 75 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 d_in[38]
port 76 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 d_in[39]
port 77 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 d_in[3]
port 78 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 d_in[40]
port 79 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 d_in[41]
port 80 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 d_in[42]
port 81 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 d_in[43]
port 82 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 d_in[44]
port 83 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 d_in[45]
port 84 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 d_in[46]
port 85 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 d_in[47]
port 86 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 d_in[48]
port 87 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 d_in[49]
port 88 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 d_in[4]
port 89 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 d_in[50]
port 90 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 d_in[51]
port 91 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 d_in[52]
port 92 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 d_in[53]
port 93 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 d_in[54]
port 94 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 d_in[55]
port 95 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 d_in[56]
port 96 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 d_in[57]
port 97 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 d_in[58]
port 98 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 d_in[59]
port 99 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 d_in[5]
port 100 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 d_in[60]
port 101 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 d_in[61]
port 102 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 d_in[62]
port 103 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 d_in[63]
port 104 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 d_in[64]
port 105 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 d_in[65]
port 106 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 d_in[66]
port 107 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 d_in[67]
port 108 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 d_in[68]
port 109 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 d_in[69]
port 110 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 d_in[6]
port 111 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 d_in[70]
port 112 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 d_in[71]
port 113 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 d_in[72]
port 114 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 d_in[73]
port 115 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 d_in[74]
port 116 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 d_in[75]
port 117 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 d_in[76]
port 118 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 d_in[77]
port 119 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 d_in[78]
port 120 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 d_in[79]
port 121 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 d_in[7]
port 122 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 d_in[80]
port 123 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 d_in[81]
port 124 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 d_in[82]
port 125 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 d_in[83]
port 126 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 d_in[84]
port 127 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 d_in[85]
port 128 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 d_in[86]
port 129 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 d_in[87]
port 130 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 d_in[88]
port 131 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 d_in[89]
port 132 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 d_in[8]
port 133 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 d_in[90]
port 134 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 d_in[91]
port 135 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 d_in[92]
port 136 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 d_in[93]
port 137 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 d_in[94]
port 138 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 d_in[95]
port 139 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 d_in[96]
port 140 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 d_in[97]
port 141 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 d_in[98]
port 142 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 d_in[99]
port 143 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 d_in[9]
port 144 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 d_out[0]
port 145 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 d_out[10]
port 146 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 d_out[11]
port 147 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 d_out[12]
port 148 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 d_out[13]
port 149 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 d_out[14]
port 150 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 d_out[15]
port 151 nsew signal output
rlabel metal2 s 113454 0 113510 800 6 d_out[16]
port 152 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 d_out[17]
port 153 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 d_out[18]
port 154 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 d_out[19]
port 155 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 d_out[1]
port 156 nsew signal output
rlabel metal2 s 116214 0 116270 800 6 d_out[20]
port 157 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 d_out[21]
port 158 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 d_out[22]
port 159 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 d_out[23]
port 160 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 d_out[24]
port 161 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 d_out[25]
port 162 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 d_out[26]
port 163 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 d_out[27]
port 164 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 d_out[28]
port 165 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 d_out[29]
port 166 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 d_out[2]
port 167 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 d_out[30]
port 168 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 d_out[31]
port 169 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 d_out[32]
port 170 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 d_out[33]
port 171 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 d_out[34]
port 172 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 d_out[35]
port 173 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 d_out[36]
port 174 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 d_out[37]
port 175 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 d_out[38]
port 176 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 d_out[39]
port 177 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 d_out[3]
port 178 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 d_out[40]
port 179 nsew signal output
rlabel metal2 s 131118 0 131174 800 6 d_out[41]
port 180 nsew signal output
rlabel metal2 s 131854 0 131910 800 6 d_out[42]
port 181 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 d_out[43]
port 182 nsew signal output
rlabel metal2 s 133234 0 133290 800 6 d_out[44]
port 183 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 d_out[45]
port 184 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 d_out[46]
port 185 nsew signal output
rlabel metal2 s 135350 0 135406 800 6 d_out[47]
port 186 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 d_out[48]
port 187 nsew signal output
rlabel metal2 s 136730 0 136786 800 6 d_out[49]
port 188 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 d_out[4]
port 189 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 d_out[50]
port 190 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 d_out[51]
port 191 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 d_out[52]
port 192 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 d_out[53]
port 193 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 d_out[54]
port 194 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 d_out[55]
port 195 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 d_out[56]
port 196 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 d_out[57]
port 197 nsew signal output
rlabel metal2 s 143170 0 143226 800 6 d_out[58]
port 198 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 d_out[59]
port 199 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 d_out[5]
port 200 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 d_out[60]
port 201 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 d_out[61]
port 202 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 d_out[62]
port 203 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 d_out[63]
port 204 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 d_out[64]
port 205 nsew signal output
rlabel metal2 s 148046 0 148102 800 6 d_out[65]
port 206 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 d_out[66]
port 207 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 d_out[67]
port 208 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 d_out[6]
port 209 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 d_out[7]
port 210 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 d_out[8]
port 211 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 d_out[9]
port 212 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 m_in[0]
port 213 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 m_in[100]
port 214 nsew signal input
rlabel metal3 s 0 77120 800 77240 6 m_in[101]
port 215 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 m_in[102]
port 216 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 m_in[103]
port 217 nsew signal input
rlabel metal3 s 0 79296 800 79416 6 m_in[104]
port 218 nsew signal input
rlabel metal3 s 0 80112 800 80232 6 m_in[105]
port 219 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 m_in[106]
port 220 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 m_in[107]
port 221 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 m_in[108]
port 222 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 m_in[109]
port 223 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 m_in[10]
port 224 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 m_in[110]
port 225 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 m_in[111]
port 226 nsew signal input
rlabel metal3 s 0 85280 800 85400 6 m_in[112]
port 227 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 m_in[113]
port 228 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 m_in[114]
port 229 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 m_in[115]
port 230 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 m_in[116]
port 231 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 m_in[117]
port 232 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 m_in[118]
port 233 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 m_in[119]
port 234 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 m_in[11]
port 235 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 m_in[120]
port 236 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 m_in[121]
port 237 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 m_in[122]
port 238 nsew signal input
rlabel metal3 s 0 93440 800 93560 6 m_in[123]
port 239 nsew signal input
rlabel metal3 s 0 94256 800 94376 6 m_in[124]
port 240 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 m_in[125]
port 241 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 m_in[126]
port 242 nsew signal input
rlabel metal3 s 0 96432 800 96552 6 m_in[127]
port 243 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 m_in[128]
port 244 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 m_in[129]
port 245 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 m_in[12]
port 246 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 m_in[130]
port 247 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 m_in[131]
port 248 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 m_in[13]
port 249 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 m_in[14]
port 250 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 m_in[15]
port 251 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 m_in[16]
port 252 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 m_in[17]
port 253 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 m_in[18]
port 254 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 m_in[19]
port 255 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 m_in[1]
port 256 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 m_in[20]
port 257 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 m_in[21]
port 258 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 m_in[22]
port 259 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 m_in[23]
port 260 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 m_in[24]
port 261 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 m_in[25]
port 262 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 m_in[26]
port 263 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 m_in[27]
port 264 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 m_in[28]
port 265 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 m_in[29]
port 266 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 m_in[2]
port 267 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 m_in[30]
port 268 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 m_in[31]
port 269 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 m_in[32]
port 270 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 m_in[33]
port 271 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 m_in[34]
port 272 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 m_in[35]
port 273 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 m_in[36]
port 274 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 m_in[37]
port 275 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 m_in[38]
port 276 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 m_in[39]
port 277 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 m_in[3]
port 278 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 m_in[40]
port 279 nsew signal input
rlabel metal3 s 0 32240 800 32360 6 m_in[41]
port 280 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 m_in[42]
port 281 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 m_in[43]
port 282 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 m_in[44]
port 283 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 m_in[45]
port 284 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 m_in[46]
port 285 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 m_in[47]
port 286 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 m_in[48]
port 287 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 m_in[49]
port 288 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 m_in[4]
port 289 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 m_in[50]
port 290 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 m_in[51]
port 291 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 m_in[52]
port 292 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 m_in[53]
port 293 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 m_in[54]
port 294 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 m_in[55]
port 295 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 m_in[56]
port 296 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 m_in[57]
port 297 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 m_in[58]
port 298 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 m_in[59]
port 299 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 m_in[5]
port 300 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 m_in[60]
port 301 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 m_in[61]
port 302 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 m_in[62]
port 303 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 m_in[63]
port 304 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 m_in[64]
port 305 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 m_in[65]
port 306 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 m_in[66]
port 307 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 m_in[67]
port 308 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 m_in[68]
port 309 nsew signal input
rlabel metal3 s 0 53184 800 53304 6 m_in[69]
port 310 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 m_in[6]
port 311 nsew signal input
rlabel metal3 s 0 54000 800 54120 6 m_in[70]
port 312 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 m_in[71]
port 313 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 m_in[72]
port 314 nsew signal input
rlabel metal3 s 0 56176 800 56296 6 m_in[73]
port 315 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 m_in[74]
port 316 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 m_in[75]
port 317 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 m_in[76]
port 318 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 m_in[77]
port 319 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 m_in[78]
port 320 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 m_in[79]
port 321 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 m_in[7]
port 322 nsew signal input
rlabel metal3 s 0 61344 800 61464 6 m_in[80]
port 323 nsew signal input
rlabel metal3 s 0 62160 800 62280 6 m_in[81]
port 324 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 m_in[82]
port 325 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 m_in[83]
port 326 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 m_in[84]
port 327 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 m_in[85]
port 328 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 m_in[86]
port 329 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 m_in[87]
port 330 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 m_in[88]
port 331 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 m_in[89]
port 332 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 m_in[8]
port 333 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 m_in[90]
port 334 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 m_in[91]
port 335 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 m_in[92]
port 336 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 m_in[93]
port 337 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 m_in[94]
port 338 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 m_in[95]
port 339 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 m_in[96]
port 340 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 m_in[97]
port 341 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 m_in[98]
port 342 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 m_in[99]
port 343 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 m_in[9]
port 344 nsew signal input
rlabel metal3 s 0 100240 800 100360 6 m_out[0]
port 345 nsew signal output
rlabel metal3 s 0 107720 800 107840 6 m_out[10]
port 346 nsew signal output
rlabel metal3 s 0 108400 800 108520 6 m_out[11]
port 347 nsew signal output
rlabel metal3 s 0 109216 800 109336 6 m_out[12]
port 348 nsew signal output
rlabel metal3 s 0 109896 800 110016 6 m_out[13]
port 349 nsew signal output
rlabel metal3 s 0 110712 800 110832 6 m_out[14]
port 350 nsew signal output
rlabel metal3 s 0 111392 800 111512 6 m_out[15]
port 351 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 m_out[16]
port 352 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 m_out[17]
port 353 nsew signal output
rlabel metal3 s 0 113704 800 113824 6 m_out[18]
port 354 nsew signal output
rlabel metal3 s 0 114384 800 114504 6 m_out[19]
port 355 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 m_out[1]
port 356 nsew signal output
rlabel metal3 s 0 115200 800 115320 6 m_out[20]
port 357 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 m_out[21]
port 358 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 m_out[22]
port 359 nsew signal output
rlabel metal3 s 0 117376 800 117496 6 m_out[23]
port 360 nsew signal output
rlabel metal3 s 0 118192 800 118312 6 m_out[24]
port 361 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 m_out[25]
port 362 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 m_out[26]
port 363 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 m_out[27]
port 364 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 m_out[28]
port 365 nsew signal output
rlabel metal3 s 0 121864 800 121984 6 m_out[29]
port 366 nsew signal output
rlabel metal3 s 0 101736 800 101856 6 m_out[2]
port 367 nsew signal output
rlabel metal3 s 0 122544 800 122664 6 m_out[30]
port 368 nsew signal output
rlabel metal3 s 0 123360 800 123480 6 m_out[31]
port 369 nsew signal output
rlabel metal3 s 0 124040 800 124160 6 m_out[32]
port 370 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 m_out[33]
port 371 nsew signal output
rlabel metal3 s 0 125536 800 125656 6 m_out[34]
port 372 nsew signal output
rlabel metal3 s 0 126352 800 126472 6 m_out[35]
port 373 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 m_out[36]
port 374 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 m_out[37]
port 375 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 m_out[38]
port 376 nsew signal output
rlabel metal3 s 0 129344 800 129464 6 m_out[39]
port 377 nsew signal output
rlabel metal3 s 0 102416 800 102536 6 m_out[3]
port 378 nsew signal output
rlabel metal3 s 0 130024 800 130144 6 m_out[40]
port 379 nsew signal output
rlabel metal3 s 0 130840 800 130960 6 m_out[41]
port 380 nsew signal output
rlabel metal3 s 0 131520 800 131640 6 m_out[42]
port 381 nsew signal output
rlabel metal3 s 0 132336 800 132456 6 m_out[43]
port 382 nsew signal output
rlabel metal3 s 0 133016 800 133136 6 m_out[44]
port 383 nsew signal output
rlabel metal3 s 0 133832 800 133952 6 m_out[45]
port 384 nsew signal output
rlabel metal3 s 0 134512 800 134632 6 m_out[46]
port 385 nsew signal output
rlabel metal3 s 0 135328 800 135448 6 m_out[47]
port 386 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 m_out[48]
port 387 nsew signal output
rlabel metal3 s 0 136824 800 136944 6 m_out[49]
port 388 nsew signal output
rlabel metal3 s 0 103232 800 103352 6 m_out[4]
port 389 nsew signal output
rlabel metal3 s 0 137504 800 137624 6 m_out[50]
port 390 nsew signal output
rlabel metal3 s 0 138320 800 138440 6 m_out[51]
port 391 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 m_out[52]
port 392 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 m_out[53]
port 393 nsew signal output
rlabel metal3 s 0 140496 800 140616 6 m_out[54]
port 394 nsew signal output
rlabel metal3 s 0 141312 800 141432 6 m_out[55]
port 395 nsew signal output
rlabel metal3 s 0 141992 800 142112 6 m_out[56]
port 396 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 m_out[57]
port 397 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 m_out[58]
port 398 nsew signal output
rlabel metal3 s 0 144304 800 144424 6 m_out[59]
port 399 nsew signal output
rlabel metal3 s 0 103912 800 104032 6 m_out[5]
port 400 nsew signal output
rlabel metal3 s 0 144984 800 145104 6 m_out[60]
port 401 nsew signal output
rlabel metal3 s 0 145800 800 145920 6 m_out[61]
port 402 nsew signal output
rlabel metal3 s 0 146480 800 146600 6 m_out[62]
port 403 nsew signal output
rlabel metal3 s 0 147296 800 147416 6 m_out[63]
port 404 nsew signal output
rlabel metal3 s 0 147976 800 148096 6 m_out[64]
port 405 nsew signal output
rlabel metal3 s 0 148792 800 148912 6 m_out[65]
port 406 nsew signal output
rlabel metal3 s 0 149472 800 149592 6 m_out[66]
port 407 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 m_out[6]
port 408 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 m_out[7]
port 409 nsew signal output
rlabel metal3 s 0 106224 800 106344 6 m_out[8]
port 410 nsew signal output
rlabel metal3 s 0 106904 800 107024 6 m_out[9]
port 411 nsew signal output
rlabel metal3 s 0 960 800 1080 6 rst
port 412 nsew signal input
rlabel metal2 s 294 0 350 800 6 stall_out
port 413 nsew signal output
rlabel metal2 s 386 149200 442 150000 6 wishbone_in[0]
port 414 nsew signal input
rlabel metal2 s 9034 149200 9090 150000 6 wishbone_in[10]
port 415 nsew signal input
rlabel metal2 s 9862 149200 9918 150000 6 wishbone_in[11]
port 416 nsew signal input
rlabel metal2 s 10782 149200 10838 150000 6 wishbone_in[12]
port 417 nsew signal input
rlabel metal2 s 11610 149200 11666 150000 6 wishbone_in[13]
port 418 nsew signal input
rlabel metal2 s 12438 149200 12494 150000 6 wishbone_in[14]
port 419 nsew signal input
rlabel metal2 s 13358 149200 13414 150000 6 wishbone_in[15]
port 420 nsew signal input
rlabel metal2 s 14186 149200 14242 150000 6 wishbone_in[16]
port 421 nsew signal input
rlabel metal2 s 15106 149200 15162 150000 6 wishbone_in[17]
port 422 nsew signal input
rlabel metal2 s 15934 149200 15990 150000 6 wishbone_in[18]
port 423 nsew signal input
rlabel metal2 s 16854 149200 16910 150000 6 wishbone_in[19]
port 424 nsew signal input
rlabel metal2 s 1214 149200 1270 150000 6 wishbone_in[1]
port 425 nsew signal input
rlabel metal2 s 17682 149200 17738 150000 6 wishbone_in[20]
port 426 nsew signal input
rlabel metal2 s 18510 149200 18566 150000 6 wishbone_in[21]
port 427 nsew signal input
rlabel metal2 s 19430 149200 19486 150000 6 wishbone_in[22]
port 428 nsew signal input
rlabel metal2 s 20258 149200 20314 150000 6 wishbone_in[23]
port 429 nsew signal input
rlabel metal2 s 21178 149200 21234 150000 6 wishbone_in[24]
port 430 nsew signal input
rlabel metal2 s 22006 149200 22062 150000 6 wishbone_in[25]
port 431 nsew signal input
rlabel metal2 s 22834 149200 22890 150000 6 wishbone_in[26]
port 432 nsew signal input
rlabel metal2 s 23754 149200 23810 150000 6 wishbone_in[27]
port 433 nsew signal input
rlabel metal2 s 24582 149200 24638 150000 6 wishbone_in[28]
port 434 nsew signal input
rlabel metal2 s 25502 149200 25558 150000 6 wishbone_in[29]
port 435 nsew signal input
rlabel metal2 s 2042 149200 2098 150000 6 wishbone_in[2]
port 436 nsew signal input
rlabel metal2 s 26330 149200 26386 150000 6 wishbone_in[30]
port 437 nsew signal input
rlabel metal2 s 27250 149200 27306 150000 6 wishbone_in[31]
port 438 nsew signal input
rlabel metal2 s 28078 149200 28134 150000 6 wishbone_in[32]
port 439 nsew signal input
rlabel metal2 s 28906 149200 28962 150000 6 wishbone_in[33]
port 440 nsew signal input
rlabel metal2 s 29826 149200 29882 150000 6 wishbone_in[34]
port 441 nsew signal input
rlabel metal2 s 30654 149200 30710 150000 6 wishbone_in[35]
port 442 nsew signal input
rlabel metal2 s 31574 149200 31630 150000 6 wishbone_in[36]
port 443 nsew signal input
rlabel metal2 s 32402 149200 32458 150000 6 wishbone_in[37]
port 444 nsew signal input
rlabel metal2 s 33322 149200 33378 150000 6 wishbone_in[38]
port 445 nsew signal input
rlabel metal2 s 34150 149200 34206 150000 6 wishbone_in[39]
port 446 nsew signal input
rlabel metal2 s 2962 149200 3018 150000 6 wishbone_in[3]
port 447 nsew signal input
rlabel metal2 s 34978 149200 35034 150000 6 wishbone_in[40]
port 448 nsew signal input
rlabel metal2 s 35898 149200 35954 150000 6 wishbone_in[41]
port 449 nsew signal input
rlabel metal2 s 36726 149200 36782 150000 6 wishbone_in[42]
port 450 nsew signal input
rlabel metal2 s 37646 149200 37702 150000 6 wishbone_in[43]
port 451 nsew signal input
rlabel metal2 s 38474 149200 38530 150000 6 wishbone_in[44]
port 452 nsew signal input
rlabel metal2 s 39302 149200 39358 150000 6 wishbone_in[45]
port 453 nsew signal input
rlabel metal2 s 40222 149200 40278 150000 6 wishbone_in[46]
port 454 nsew signal input
rlabel metal2 s 41050 149200 41106 150000 6 wishbone_in[47]
port 455 nsew signal input
rlabel metal2 s 41970 149200 42026 150000 6 wishbone_in[48]
port 456 nsew signal input
rlabel metal2 s 42798 149200 42854 150000 6 wishbone_in[49]
port 457 nsew signal input
rlabel metal2 s 3790 149200 3846 150000 6 wishbone_in[4]
port 458 nsew signal input
rlabel metal2 s 43718 149200 43774 150000 6 wishbone_in[50]
port 459 nsew signal input
rlabel metal2 s 44546 149200 44602 150000 6 wishbone_in[51]
port 460 nsew signal input
rlabel metal2 s 45374 149200 45430 150000 6 wishbone_in[52]
port 461 nsew signal input
rlabel metal2 s 46294 149200 46350 150000 6 wishbone_in[53]
port 462 nsew signal input
rlabel metal2 s 47122 149200 47178 150000 6 wishbone_in[54]
port 463 nsew signal input
rlabel metal2 s 48042 149200 48098 150000 6 wishbone_in[55]
port 464 nsew signal input
rlabel metal2 s 48870 149200 48926 150000 6 wishbone_in[56]
port 465 nsew signal input
rlabel metal2 s 49790 149200 49846 150000 6 wishbone_in[57]
port 466 nsew signal input
rlabel metal2 s 50618 149200 50674 150000 6 wishbone_in[58]
port 467 nsew signal input
rlabel metal2 s 51446 149200 51502 150000 6 wishbone_in[59]
port 468 nsew signal input
rlabel metal2 s 4710 149200 4766 150000 6 wishbone_in[5]
port 469 nsew signal input
rlabel metal2 s 52366 149200 52422 150000 6 wishbone_in[60]
port 470 nsew signal input
rlabel metal2 s 53194 149200 53250 150000 6 wishbone_in[61]
port 471 nsew signal input
rlabel metal2 s 54114 149200 54170 150000 6 wishbone_in[62]
port 472 nsew signal input
rlabel metal2 s 54942 149200 54998 150000 6 wishbone_in[63]
port 473 nsew signal input
rlabel metal2 s 55862 149200 55918 150000 6 wishbone_in[64]
port 474 nsew signal input
rlabel metal2 s 56690 149200 56746 150000 6 wishbone_in[65]
port 475 nsew signal input
rlabel metal2 s 5538 149200 5594 150000 6 wishbone_in[6]
port 476 nsew signal input
rlabel metal2 s 6366 149200 6422 150000 6 wishbone_in[7]
port 477 nsew signal input
rlabel metal2 s 7286 149200 7342 150000 6 wishbone_in[8]
port 478 nsew signal input
rlabel metal2 s 8114 149200 8170 150000 6 wishbone_in[9]
port 479 nsew signal input
rlabel metal2 s 57518 149200 57574 150000 6 wishbone_out[0]
port 480 nsew signal output
rlabel metal2 s 144274 149200 144330 150000 6 wishbone_out[100]
port 481 nsew signal output
rlabel metal2 s 145102 149200 145158 150000 6 wishbone_out[101]
port 482 nsew signal output
rlabel metal2 s 145930 149200 145986 150000 6 wishbone_out[102]
port 483 nsew signal output
rlabel metal2 s 146850 149200 146906 150000 6 wishbone_out[103]
port 484 nsew signal output
rlabel metal2 s 147678 149200 147734 150000 6 wishbone_out[104]
port 485 nsew signal output
rlabel metal2 s 148598 149200 148654 150000 6 wishbone_out[105]
port 486 nsew signal output
rlabel metal2 s 149426 149200 149482 150000 6 wishbone_out[106]
port 487 nsew signal output
rlabel metal2 s 66258 149200 66314 150000 6 wishbone_out[10]
port 488 nsew signal output
rlabel metal2 s 67086 149200 67142 150000 6 wishbone_out[11]
port 489 nsew signal output
rlabel metal2 s 67914 149200 67970 150000 6 wishbone_out[12]
port 490 nsew signal output
rlabel metal2 s 68834 149200 68890 150000 6 wishbone_out[13]
port 491 nsew signal output
rlabel metal2 s 69662 149200 69718 150000 6 wishbone_out[14]
port 492 nsew signal output
rlabel metal2 s 70582 149200 70638 150000 6 wishbone_out[15]
port 493 nsew signal output
rlabel metal2 s 71410 149200 71466 150000 6 wishbone_out[16]
port 494 nsew signal output
rlabel metal2 s 72330 149200 72386 150000 6 wishbone_out[17]
port 495 nsew signal output
rlabel metal2 s 73158 149200 73214 150000 6 wishbone_out[18]
port 496 nsew signal output
rlabel metal2 s 73986 149200 74042 150000 6 wishbone_out[19]
port 497 nsew signal output
rlabel metal2 s 58438 149200 58494 150000 6 wishbone_out[1]
port 498 nsew signal output
rlabel metal2 s 74906 149200 74962 150000 6 wishbone_out[20]
port 499 nsew signal output
rlabel metal2 s 75734 149200 75790 150000 6 wishbone_out[21]
port 500 nsew signal output
rlabel metal2 s 76654 149200 76710 150000 6 wishbone_out[22]
port 501 nsew signal output
rlabel metal2 s 77482 149200 77538 150000 6 wishbone_out[23]
port 502 nsew signal output
rlabel metal2 s 78310 149200 78366 150000 6 wishbone_out[24]
port 503 nsew signal output
rlabel metal2 s 79230 149200 79286 150000 6 wishbone_out[25]
port 504 nsew signal output
rlabel metal2 s 80058 149200 80114 150000 6 wishbone_out[26]
port 505 nsew signal output
rlabel metal2 s 80978 149200 81034 150000 6 wishbone_out[27]
port 506 nsew signal output
rlabel metal2 s 81806 149200 81862 150000 6 wishbone_out[28]
port 507 nsew signal output
rlabel metal2 s 82726 149200 82782 150000 6 wishbone_out[29]
port 508 nsew signal output
rlabel metal2 s 59266 149200 59322 150000 6 wishbone_out[2]
port 509 nsew signal output
rlabel metal2 s 83554 149200 83610 150000 6 wishbone_out[30]
port 510 nsew signal output
rlabel metal2 s 84382 149200 84438 150000 6 wishbone_out[31]
port 511 nsew signal output
rlabel metal2 s 85302 149200 85358 150000 6 wishbone_out[32]
port 512 nsew signal output
rlabel metal2 s 86130 149200 86186 150000 6 wishbone_out[33]
port 513 nsew signal output
rlabel metal2 s 87050 149200 87106 150000 6 wishbone_out[34]
port 514 nsew signal output
rlabel metal2 s 87878 149200 87934 150000 6 wishbone_out[35]
port 515 nsew signal output
rlabel metal2 s 88798 149200 88854 150000 6 wishbone_out[36]
port 516 nsew signal output
rlabel metal2 s 89626 149200 89682 150000 6 wishbone_out[37]
port 517 nsew signal output
rlabel metal2 s 90454 149200 90510 150000 6 wishbone_out[38]
port 518 nsew signal output
rlabel metal2 s 91374 149200 91430 150000 6 wishbone_out[39]
port 519 nsew signal output
rlabel metal2 s 60186 149200 60242 150000 6 wishbone_out[3]
port 520 nsew signal output
rlabel metal2 s 92202 149200 92258 150000 6 wishbone_out[40]
port 521 nsew signal output
rlabel metal2 s 93122 149200 93178 150000 6 wishbone_out[41]
port 522 nsew signal output
rlabel metal2 s 93950 149200 94006 150000 6 wishbone_out[42]
port 523 nsew signal output
rlabel metal2 s 94778 149200 94834 150000 6 wishbone_out[43]
port 524 nsew signal output
rlabel metal2 s 95698 149200 95754 150000 6 wishbone_out[44]
port 525 nsew signal output
rlabel metal2 s 96526 149200 96582 150000 6 wishbone_out[45]
port 526 nsew signal output
rlabel metal2 s 97446 149200 97502 150000 6 wishbone_out[46]
port 527 nsew signal output
rlabel metal2 s 98274 149200 98330 150000 6 wishbone_out[47]
port 528 nsew signal output
rlabel metal2 s 99194 149200 99250 150000 6 wishbone_out[48]
port 529 nsew signal output
rlabel metal2 s 100022 149200 100078 150000 6 wishbone_out[49]
port 530 nsew signal output
rlabel metal2 s 61014 149200 61070 150000 6 wishbone_out[4]
port 531 nsew signal output
rlabel metal2 s 100850 149200 100906 150000 6 wishbone_out[50]
port 532 nsew signal output
rlabel metal2 s 101770 149200 101826 150000 6 wishbone_out[51]
port 533 nsew signal output
rlabel metal2 s 102598 149200 102654 150000 6 wishbone_out[52]
port 534 nsew signal output
rlabel metal2 s 103518 149200 103574 150000 6 wishbone_out[53]
port 535 nsew signal output
rlabel metal2 s 104346 149200 104402 150000 6 wishbone_out[54]
port 536 nsew signal output
rlabel metal2 s 105266 149200 105322 150000 6 wishbone_out[55]
port 537 nsew signal output
rlabel metal2 s 106094 149200 106150 150000 6 wishbone_out[56]
port 538 nsew signal output
rlabel metal2 s 106922 149200 106978 150000 6 wishbone_out[57]
port 539 nsew signal output
rlabel metal2 s 107842 149200 107898 150000 6 wishbone_out[58]
port 540 nsew signal output
rlabel metal2 s 108670 149200 108726 150000 6 wishbone_out[59]
port 541 nsew signal output
rlabel metal2 s 61842 149200 61898 150000 6 wishbone_out[5]
port 542 nsew signal output
rlabel metal2 s 109590 149200 109646 150000 6 wishbone_out[60]
port 543 nsew signal output
rlabel metal2 s 110418 149200 110474 150000 6 wishbone_out[61]
port 544 nsew signal output
rlabel metal2 s 111338 149200 111394 150000 6 wishbone_out[62]
port 545 nsew signal output
rlabel metal2 s 112166 149200 112222 150000 6 wishbone_out[63]
port 546 nsew signal output
rlabel metal2 s 112994 149200 113050 150000 6 wishbone_out[64]
port 547 nsew signal output
rlabel metal2 s 113914 149200 113970 150000 6 wishbone_out[65]
port 548 nsew signal output
rlabel metal2 s 114742 149200 114798 150000 6 wishbone_out[66]
port 549 nsew signal output
rlabel metal2 s 115662 149200 115718 150000 6 wishbone_out[67]
port 550 nsew signal output
rlabel metal2 s 116490 149200 116546 150000 6 wishbone_out[68]
port 551 nsew signal output
rlabel metal2 s 117318 149200 117374 150000 6 wishbone_out[69]
port 552 nsew signal output
rlabel metal2 s 62762 149200 62818 150000 6 wishbone_out[6]
port 553 nsew signal output
rlabel metal2 s 118238 149200 118294 150000 6 wishbone_out[70]
port 554 nsew signal output
rlabel metal2 s 119066 149200 119122 150000 6 wishbone_out[71]
port 555 nsew signal output
rlabel metal2 s 119986 149200 120042 150000 6 wishbone_out[72]
port 556 nsew signal output
rlabel metal2 s 120814 149200 120870 150000 6 wishbone_out[73]
port 557 nsew signal output
rlabel metal2 s 121734 149200 121790 150000 6 wishbone_out[74]
port 558 nsew signal output
rlabel metal2 s 122562 149200 122618 150000 6 wishbone_out[75]
port 559 nsew signal output
rlabel metal2 s 123390 149200 123446 150000 6 wishbone_out[76]
port 560 nsew signal output
rlabel metal2 s 124310 149200 124366 150000 6 wishbone_out[77]
port 561 nsew signal output
rlabel metal2 s 125138 149200 125194 150000 6 wishbone_out[78]
port 562 nsew signal output
rlabel metal2 s 126058 149200 126114 150000 6 wishbone_out[79]
port 563 nsew signal output
rlabel metal2 s 63590 149200 63646 150000 6 wishbone_out[7]
port 564 nsew signal output
rlabel metal2 s 126886 149200 126942 150000 6 wishbone_out[80]
port 565 nsew signal output
rlabel metal2 s 127806 149200 127862 150000 6 wishbone_out[81]
port 566 nsew signal output
rlabel metal2 s 128634 149200 128690 150000 6 wishbone_out[82]
port 567 nsew signal output
rlabel metal2 s 129462 149200 129518 150000 6 wishbone_out[83]
port 568 nsew signal output
rlabel metal2 s 130382 149200 130438 150000 6 wishbone_out[84]
port 569 nsew signal output
rlabel metal2 s 131210 149200 131266 150000 6 wishbone_out[85]
port 570 nsew signal output
rlabel metal2 s 132130 149200 132186 150000 6 wishbone_out[86]
port 571 nsew signal output
rlabel metal2 s 132958 149200 133014 150000 6 wishbone_out[87]
port 572 nsew signal output
rlabel metal2 s 133786 149200 133842 150000 6 wishbone_out[88]
port 573 nsew signal output
rlabel metal2 s 134706 149200 134762 150000 6 wishbone_out[89]
port 574 nsew signal output
rlabel metal2 s 64510 149200 64566 150000 6 wishbone_out[8]
port 575 nsew signal output
rlabel metal2 s 135534 149200 135590 150000 6 wishbone_out[90]
port 576 nsew signal output
rlabel metal2 s 136454 149200 136510 150000 6 wishbone_out[91]
port 577 nsew signal output
rlabel metal2 s 137282 149200 137338 150000 6 wishbone_out[92]
port 578 nsew signal output
rlabel metal2 s 138202 149200 138258 150000 6 wishbone_out[93]
port 579 nsew signal output
rlabel metal2 s 139030 149200 139086 150000 6 wishbone_out[94]
port 580 nsew signal output
rlabel metal2 s 139858 149200 139914 150000 6 wishbone_out[95]
port 581 nsew signal output
rlabel metal2 s 140778 149200 140834 150000 6 wishbone_out[96]
port 582 nsew signal output
rlabel metal2 s 141606 149200 141662 150000 6 wishbone_out[97]
port 583 nsew signal output
rlabel metal2 s 142526 149200 142582 150000 6 wishbone_out[98]
port 584 nsew signal output
rlabel metal2 s 143354 149200 143410 150000 6 wishbone_out[99]
port 585 nsew signal output
rlabel metal2 s 65338 149200 65394 150000 6 wishbone_out[9]
port 586 nsew signal output
rlabel metal4 s 127088 2128 127408 147472 6 vccd1
port 587 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 147472 6 vccd1
port 588 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 147472 6 vccd1
port 589 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 147472 6 vccd1
port 590 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 147472 6 vccd1
port 591 nsew power bidirectional
rlabel metal4 s 142448 2128 142768 147472 6 vssd1
port 592 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 147472 6 vssd1
port 593 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 147472 6 vssd1
port 594 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 147472 6 vssd1
port 595 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 147472 6 vssd1
port 596 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 150000 150000
string LEFview TRUE
string GDS_FILE /project/openlane/dcache/runs/dcache/results/magic/dcache.gds
string GDS_END 69473548
string GDS_START 406954
<< end >>

