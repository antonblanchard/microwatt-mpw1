VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiply_4
  CLASS BLOCK ;
  FOREIGN multiply_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 1100.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 1096.000 2.210 1100.000 ;
    END
  END clk
  PIN m_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 1096.000 6.350 1100.000 ;
    END
  END m_in[0]
  PIN m_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 1096.000 429.090 1100.000 ;
    END
  END m_in[100]
  PIN m_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 1096.000 433.690 1100.000 ;
    END
  END m_in[101]
  PIN m_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 1096.000 437.830 1100.000 ;
    END
  END m_in[102]
  PIN m_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 1096.000 441.970 1100.000 ;
    END
  END m_in[103]
  PIN m_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 1096.000 446.110 1100.000 ;
    END
  END m_in[104]
  PIN m_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 1096.000 450.250 1100.000 ;
    END
  END m_in[105]
  PIN m_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1096.000 454.390 1100.000 ;
    END
  END m_in[106]
  PIN m_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 1096.000 458.990 1100.000 ;
    END
  END m_in[107]
  PIN m_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 1096.000 463.130 1100.000 ;
    END
  END m_in[108]
  PIN m_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 1096.000 467.270 1100.000 ;
    END
  END m_in[109]
  PIN m_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1096.000 48.670 1100.000 ;
    END
  END m_in[10]
  PIN m_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 1096.000 471.410 1100.000 ;
    END
  END m_in[110]
  PIN m_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 1096.000 475.550 1100.000 ;
    END
  END m_in[111]
  PIN m_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1096.000 480.150 1100.000 ;
    END
  END m_in[112]
  PIN m_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 1096.000 484.290 1100.000 ;
    END
  END m_in[113]
  PIN m_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 1096.000 488.430 1100.000 ;
    END
  END m_in[114]
  PIN m_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 1096.000 492.570 1100.000 ;
    END
  END m_in[115]
  PIN m_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 1096.000 496.710 1100.000 ;
    END
  END m_in[116]
  PIN m_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 1096.000 501.310 1100.000 ;
    END
  END m_in[117]
  PIN m_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 1096.000 505.450 1100.000 ;
    END
  END m_in[118]
  PIN m_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 1096.000 509.590 1100.000 ;
    END
  END m_in[119]
  PIN m_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 1096.000 52.810 1100.000 ;
    END
  END m_in[11]
  PIN m_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 1096.000 513.730 1100.000 ;
    END
  END m_in[120]
  PIN m_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 1096.000 517.870 1100.000 ;
    END
  END m_in[121]
  PIN m_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 1096.000 522.470 1100.000 ;
    END
  END m_in[122]
  PIN m_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 1096.000 526.610 1100.000 ;
    END
  END m_in[123]
  PIN m_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 1096.000 530.750 1100.000 ;
    END
  END m_in[124]
  PIN m_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 1096.000 534.890 1100.000 ;
    END
  END m_in[125]
  PIN m_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 1096.000 539.030 1100.000 ;
    END
  END m_in[126]
  PIN m_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 1096.000 543.630 1100.000 ;
    END
  END m_in[127]
  PIN m_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 1096.000 547.770 1100.000 ;
    END
  END m_in[128]
  PIN m_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 1096.000 551.910 1100.000 ;
    END
  END m_in[129]
  PIN m_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 1096.000 56.950 1100.000 ;
    END
  END m_in[12]
  PIN m_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 1096.000 556.050 1100.000 ;
    END
  END m_in[130]
  PIN m_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 1096.000 560.190 1100.000 ;
    END
  END m_in[131]
  PIN m_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 1096.000 564.790 1100.000 ;
    END
  END m_in[132]
  PIN m_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 1096.000 568.930 1100.000 ;
    END
  END m_in[133]
  PIN m_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 1096.000 573.070 1100.000 ;
    END
  END m_in[134]
  PIN m_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 1096.000 577.210 1100.000 ;
    END
  END m_in[135]
  PIN m_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 1096.000 581.350 1100.000 ;
    END
  END m_in[136]
  PIN m_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 1096.000 585.950 1100.000 ;
    END
  END m_in[137]
  PIN m_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 1096.000 590.090 1100.000 ;
    END
  END m_in[138]
  PIN m_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 1096.000 594.230 1100.000 ;
    END
  END m_in[139]
  PIN m_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 1096.000 61.090 1100.000 ;
    END
  END m_in[13]
  PIN m_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 1096.000 598.370 1100.000 ;
    END
  END m_in[140]
  PIN m_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 1096.000 602.510 1100.000 ;
    END
  END m_in[141]
  PIN m_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 1096.000 607.110 1100.000 ;
    END
  END m_in[142]
  PIN m_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 1096.000 611.250 1100.000 ;
    END
  END m_in[143]
  PIN m_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1096.000 615.390 1100.000 ;
    END
  END m_in[144]
  PIN m_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 1096.000 619.530 1100.000 ;
    END
  END m_in[145]
  PIN m_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 1096.000 623.670 1100.000 ;
    END
  END m_in[146]
  PIN m_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 1096.000 628.270 1100.000 ;
    END
  END m_in[147]
  PIN m_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 1096.000 632.410 1100.000 ;
    END
  END m_in[148]
  PIN m_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 1096.000 636.550 1100.000 ;
    END
  END m_in[149]
  PIN m_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 1096.000 65.230 1100.000 ;
    END
  END m_in[14]
  PIN m_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 1096.000 640.690 1100.000 ;
    END
  END m_in[150]
  PIN m_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 1096.000 644.830 1100.000 ;
    END
  END m_in[151]
  PIN m_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 1096.000 649.430 1100.000 ;
    END
  END m_in[152]
  PIN m_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 1096.000 653.570 1100.000 ;
    END
  END m_in[153]
  PIN m_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 1096.000 657.710 1100.000 ;
    END
  END m_in[154]
  PIN m_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 1096.000 661.850 1100.000 ;
    END
  END m_in[155]
  PIN m_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 1096.000 665.990 1100.000 ;
    END
  END m_in[156]
  PIN m_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 1096.000 670.130 1100.000 ;
    END
  END m_in[157]
  PIN m_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 1096.000 674.730 1100.000 ;
    END
  END m_in[158]
  PIN m_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 1096.000 678.870 1100.000 ;
    END
  END m_in[159]
  PIN m_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 1096.000 69.830 1100.000 ;
    END
  END m_in[15]
  PIN m_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 1096.000 683.010 1100.000 ;
    END
  END m_in[160]
  PIN m_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 1096.000 687.150 1100.000 ;
    END
  END m_in[161]
  PIN m_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 1096.000 691.290 1100.000 ;
    END
  END m_in[162]
  PIN m_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 1096.000 695.890 1100.000 ;
    END
  END m_in[163]
  PIN m_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 1096.000 700.030 1100.000 ;
    END
  END m_in[164]
  PIN m_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 1096.000 704.170 1100.000 ;
    END
  END m_in[165]
  PIN m_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 1096.000 708.310 1100.000 ;
    END
  END m_in[166]
  PIN m_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 1096.000 712.450 1100.000 ;
    END
  END m_in[167]
  PIN m_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 1096.000 717.050 1100.000 ;
    END
  END m_in[168]
  PIN m_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 1096.000 721.190 1100.000 ;
    END
  END m_in[169]
  PIN m_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 1096.000 73.970 1100.000 ;
    END
  END m_in[16]
  PIN m_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 1096.000 725.330 1100.000 ;
    END
  END m_in[170]
  PIN m_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 1096.000 729.470 1100.000 ;
    END
  END m_in[171]
  PIN m_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 1096.000 733.610 1100.000 ;
    END
  END m_in[172]
  PIN m_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 1096.000 738.210 1100.000 ;
    END
  END m_in[173]
  PIN m_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 1096.000 742.350 1100.000 ;
    END
  END m_in[174]
  PIN m_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 1096.000 746.490 1100.000 ;
    END
  END m_in[175]
  PIN m_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 1096.000 750.630 1100.000 ;
    END
  END m_in[176]
  PIN m_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 1096.000 754.770 1100.000 ;
    END
  END m_in[177]
  PIN m_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 1096.000 759.370 1100.000 ;
    END
  END m_in[178]
  PIN m_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1096.000 763.510 1100.000 ;
    END
  END m_in[179]
  PIN m_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 1096.000 78.110 1100.000 ;
    END
  END m_in[17]
  PIN m_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 1096.000 767.650 1100.000 ;
    END
  END m_in[180]
  PIN m_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 1096.000 771.790 1100.000 ;
    END
  END m_in[181]
  PIN m_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 1096.000 775.930 1100.000 ;
    END
  END m_in[182]
  PIN m_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 1096.000 780.530 1100.000 ;
    END
  END m_in[183]
  PIN m_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 1096.000 784.670 1100.000 ;
    END
  END m_in[184]
  PIN m_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 1096.000 788.810 1100.000 ;
    END
  END m_in[185]
  PIN m_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 1096.000 792.950 1100.000 ;
    END
  END m_in[186]
  PIN m_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 1096.000 797.090 1100.000 ;
    END
  END m_in[187]
  PIN m_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 1096.000 801.690 1100.000 ;
    END
  END m_in[188]
  PIN m_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 1096.000 805.830 1100.000 ;
    END
  END m_in[189]
  PIN m_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 1096.000 82.250 1100.000 ;
    END
  END m_in[18]
  PIN m_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 1096.000 809.970 1100.000 ;
    END
  END m_in[190]
  PIN m_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 1096.000 814.110 1100.000 ;
    END
  END m_in[191]
  PIN m_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 1096.000 818.250 1100.000 ;
    END
  END m_in[192]
  PIN m_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 1096.000 822.850 1100.000 ;
    END
  END m_in[193]
  PIN m_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 1096.000 826.990 1100.000 ;
    END
  END m_in[194]
  PIN m_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 1096.000 831.130 1100.000 ;
    END
  END m_in[195]
  PIN m_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 1096.000 835.270 1100.000 ;
    END
  END m_in[196]
  PIN m_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 1096.000 839.410 1100.000 ;
    END
  END m_in[197]
  PIN m_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 1096.000 844.010 1100.000 ;
    END
  END m_in[198]
  PIN m_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.870 1096.000 848.150 1100.000 ;
    END
  END m_in[199]
  PIN m_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 1096.000 86.390 1100.000 ;
    END
  END m_in[19]
  PIN m_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 1096.000 10.490 1100.000 ;
    END
  END m_in[1]
  PIN m_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 1096.000 852.290 1100.000 ;
    END
  END m_in[200]
  PIN m_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 1096.000 856.430 1100.000 ;
    END
  END m_in[201]
  PIN m_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 1096.000 860.570 1100.000 ;
    END
  END m_in[202]
  PIN m_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 1096.000 865.170 1100.000 ;
    END
  END m_in[203]
  PIN m_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 1096.000 869.310 1100.000 ;
    END
  END m_in[204]
  PIN m_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 1096.000 873.450 1100.000 ;
    END
  END m_in[205]
  PIN m_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 1096.000 877.590 1100.000 ;
    END
  END m_in[206]
  PIN m_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 1096.000 881.730 1100.000 ;
    END
  END m_in[207]
  PIN m_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 1096.000 885.870 1100.000 ;
    END
  END m_in[208]
  PIN m_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 1096.000 890.470 1100.000 ;
    END
  END m_in[209]
  PIN m_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 1096.000 90.990 1100.000 ;
    END
  END m_in[20]
  PIN m_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 1096.000 894.610 1100.000 ;
    END
  END m_in[210]
  PIN m_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 1096.000 898.750 1100.000 ;
    END
  END m_in[211]
  PIN m_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 1096.000 902.890 1100.000 ;
    END
  END m_in[212]
  PIN m_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 1096.000 907.030 1100.000 ;
    END
  END m_in[213]
  PIN m_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 1096.000 911.630 1100.000 ;
    END
  END m_in[214]
  PIN m_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 1096.000 915.770 1100.000 ;
    END
  END m_in[215]
  PIN m_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 1096.000 919.910 1100.000 ;
    END
  END m_in[216]
  PIN m_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 1096.000 924.050 1100.000 ;
    END
  END m_in[217]
  PIN m_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 1096.000 928.190 1100.000 ;
    END
  END m_in[218]
  PIN m_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 1096.000 932.790 1100.000 ;
    END
  END m_in[219]
  PIN m_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 1096.000 95.130 1100.000 ;
    END
  END m_in[21]
  PIN m_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 1096.000 936.930 1100.000 ;
    END
  END m_in[220]
  PIN m_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.790 1096.000 941.070 1100.000 ;
    END
  END m_in[221]
  PIN m_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 1096.000 945.210 1100.000 ;
    END
  END m_in[222]
  PIN m_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 1096.000 949.350 1100.000 ;
    END
  END m_in[223]
  PIN m_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 1096.000 953.950 1100.000 ;
    END
  END m_in[224]
  PIN m_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 1096.000 958.090 1100.000 ;
    END
  END m_in[225]
  PIN m_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 1096.000 962.230 1100.000 ;
    END
  END m_in[226]
  PIN m_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 1096.000 966.370 1100.000 ;
    END
  END m_in[227]
  PIN m_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 1096.000 970.510 1100.000 ;
    END
  END m_in[228]
  PIN m_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 1096.000 975.110 1100.000 ;
    END
  END m_in[229]
  PIN m_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 1096.000 99.270 1100.000 ;
    END
  END m_in[22]
  PIN m_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 1096.000 979.250 1100.000 ;
    END
  END m_in[230]
  PIN m_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 1096.000 983.390 1100.000 ;
    END
  END m_in[231]
  PIN m_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 1096.000 987.530 1100.000 ;
    END
  END m_in[232]
  PIN m_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 1096.000 991.670 1100.000 ;
    END
  END m_in[233]
  PIN m_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 1096.000 996.270 1100.000 ;
    END
  END m_in[234]
  PIN m_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.130 1096.000 1000.410 1100.000 ;
    END
  END m_in[235]
  PIN m_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.270 1096.000 1004.550 1100.000 ;
    END
  END m_in[236]
  PIN m_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 1096.000 1008.690 1100.000 ;
    END
  END m_in[237]
  PIN m_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 1096.000 1012.830 1100.000 ;
    END
  END m_in[238]
  PIN m_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 1096.000 1017.430 1100.000 ;
    END
  END m_in[239]
  PIN m_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1096.000 103.410 1100.000 ;
    END
  END m_in[23]
  PIN m_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 1096.000 1021.570 1100.000 ;
    END
  END m_in[240]
  PIN m_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.430 1096.000 1025.710 1100.000 ;
    END
  END m_in[241]
  PIN m_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 1096.000 1029.850 1100.000 ;
    END
  END m_in[242]
  PIN m_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 1096.000 1033.990 1100.000 ;
    END
  END m_in[243]
  PIN m_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 1096.000 1038.590 1100.000 ;
    END
  END m_in[244]
  PIN m_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.450 1096.000 1042.730 1100.000 ;
    END
  END m_in[245]
  PIN m_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 1096.000 1046.870 1100.000 ;
    END
  END m_in[246]
  PIN m_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 1096.000 1051.010 1100.000 ;
    END
  END m_in[247]
  PIN m_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.870 1096.000 1055.150 1100.000 ;
    END
  END m_in[248]
  PIN m_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 1096.000 1059.750 1100.000 ;
    END
  END m_in[249]
  PIN m_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 1096.000 107.550 1100.000 ;
    END
  END m_in[24]
  PIN m_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.610 1096.000 1063.890 1100.000 ;
    END
  END m_in[250]
  PIN m_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 1096.000 1068.030 1100.000 ;
    END
  END m_in[251]
  PIN m_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 1096.000 1072.170 1100.000 ;
    END
  END m_in[252]
  PIN m_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.030 1096.000 1076.310 1100.000 ;
    END
  END m_in[253]
  PIN m_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 1096.000 1080.910 1100.000 ;
    END
  END m_in[254]
  PIN m_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.770 1096.000 1085.050 1100.000 ;
    END
  END m_in[255]
  PIN m_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 1096.000 1089.190 1100.000 ;
    END
  END m_in[256]
  PIN m_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 1096.000 1093.330 1100.000 ;
    END
  END m_in[257]
  PIN m_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.190 1096.000 1097.470 1100.000 ;
    END
  END m_in[258]
  PIN m_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 1096.000 112.150 1100.000 ;
    END
  END m_in[25]
  PIN m_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 1096.000 116.290 1100.000 ;
    END
  END m_in[26]
  PIN m_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 1096.000 120.430 1100.000 ;
    END
  END m_in[27]
  PIN m_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 1096.000 124.570 1100.000 ;
    END
  END m_in[28]
  PIN m_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 1096.000 128.710 1100.000 ;
    END
  END m_in[29]
  PIN m_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 1096.000 14.630 1100.000 ;
    END
  END m_in[2]
  PIN m_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 1096.000 133.310 1100.000 ;
    END
  END m_in[30]
  PIN m_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 1096.000 137.450 1100.000 ;
    END
  END m_in[31]
  PIN m_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 1096.000 141.590 1100.000 ;
    END
  END m_in[32]
  PIN m_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 1096.000 145.730 1100.000 ;
    END
  END m_in[33]
  PIN m_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 1096.000 149.870 1100.000 ;
    END
  END m_in[34]
  PIN m_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 1096.000 154.470 1100.000 ;
    END
  END m_in[35]
  PIN m_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 1096.000 158.610 1100.000 ;
    END
  END m_in[36]
  PIN m_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 1096.000 162.750 1100.000 ;
    END
  END m_in[37]
  PIN m_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 1096.000 166.890 1100.000 ;
    END
  END m_in[38]
  PIN m_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 1096.000 171.030 1100.000 ;
    END
  END m_in[39]
  PIN m_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 1096.000 18.770 1100.000 ;
    END
  END m_in[3]
  PIN m_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 1096.000 175.630 1100.000 ;
    END
  END m_in[40]
  PIN m_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 1096.000 179.770 1100.000 ;
    END
  END m_in[41]
  PIN m_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 1096.000 183.910 1100.000 ;
    END
  END m_in[42]
  PIN m_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 1096.000 188.050 1100.000 ;
    END
  END m_in[43]
  PIN m_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 1096.000 192.190 1100.000 ;
    END
  END m_in[44]
  PIN m_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 1096.000 196.790 1100.000 ;
    END
  END m_in[45]
  PIN m_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 1096.000 200.930 1100.000 ;
    END
  END m_in[46]
  PIN m_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 1096.000 205.070 1100.000 ;
    END
  END m_in[47]
  PIN m_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 1096.000 209.210 1100.000 ;
    END
  END m_in[48]
  PIN m_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 1096.000 213.350 1100.000 ;
    END
  END m_in[49]
  PIN m_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1096.000 22.910 1100.000 ;
    END
  END m_in[4]
  PIN m_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 1096.000 217.950 1100.000 ;
    END
  END m_in[50]
  PIN m_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 1096.000 222.090 1100.000 ;
    END
  END m_in[51]
  PIN m_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 1096.000 226.230 1100.000 ;
    END
  END m_in[52]
  PIN m_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 1096.000 230.370 1100.000 ;
    END
  END m_in[53]
  PIN m_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 1096.000 234.510 1100.000 ;
    END
  END m_in[54]
  PIN m_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 1096.000 238.650 1100.000 ;
    END
  END m_in[55]
  PIN m_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 1096.000 243.250 1100.000 ;
    END
  END m_in[56]
  PIN m_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 1096.000 247.390 1100.000 ;
    END
  END m_in[57]
  PIN m_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1096.000 251.530 1100.000 ;
    END
  END m_in[58]
  PIN m_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 1096.000 255.670 1100.000 ;
    END
  END m_in[59]
  PIN m_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 1096.000 27.510 1100.000 ;
    END
  END m_in[5]
  PIN m_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 1096.000 259.810 1100.000 ;
    END
  END m_in[60]
  PIN m_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 1096.000 264.410 1100.000 ;
    END
  END m_in[61]
  PIN m_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 1096.000 268.550 1100.000 ;
    END
  END m_in[62]
  PIN m_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 1096.000 272.690 1100.000 ;
    END
  END m_in[63]
  PIN m_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 1096.000 276.830 1100.000 ;
    END
  END m_in[64]
  PIN m_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 1096.000 280.970 1100.000 ;
    END
  END m_in[65]
  PIN m_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 1096.000 285.570 1100.000 ;
    END
  END m_in[66]
  PIN m_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 1096.000 289.710 1100.000 ;
    END
  END m_in[67]
  PIN m_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 1096.000 293.850 1100.000 ;
    END
  END m_in[68]
  PIN m_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 1096.000 297.990 1100.000 ;
    END
  END m_in[69]
  PIN m_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 1096.000 31.650 1100.000 ;
    END
  END m_in[6]
  PIN m_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 1096.000 302.130 1100.000 ;
    END
  END m_in[70]
  PIN m_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 1096.000 306.730 1100.000 ;
    END
  END m_in[71]
  PIN m_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 1096.000 310.870 1100.000 ;
    END
  END m_in[72]
  PIN m_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 1096.000 315.010 1100.000 ;
    END
  END m_in[73]
  PIN m_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 1096.000 319.150 1100.000 ;
    END
  END m_in[74]
  PIN m_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 1096.000 323.290 1100.000 ;
    END
  END m_in[75]
  PIN m_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 1096.000 327.890 1100.000 ;
    END
  END m_in[76]
  PIN m_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 1096.000 332.030 1100.000 ;
    END
  END m_in[77]
  PIN m_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 1096.000 336.170 1100.000 ;
    END
  END m_in[78]
  PIN m_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 1096.000 340.310 1100.000 ;
    END
  END m_in[79]
  PIN m_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1096.000 35.790 1100.000 ;
    END
  END m_in[7]
  PIN m_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 1096.000 344.450 1100.000 ;
    END
  END m_in[80]
  PIN m_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 1096.000 349.050 1100.000 ;
    END
  END m_in[81]
  PIN m_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 1096.000 353.190 1100.000 ;
    END
  END m_in[82]
  PIN m_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 1096.000 357.330 1100.000 ;
    END
  END m_in[83]
  PIN m_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 1096.000 361.470 1100.000 ;
    END
  END m_in[84]
  PIN m_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 1096.000 365.610 1100.000 ;
    END
  END m_in[85]
  PIN m_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 1096.000 370.210 1100.000 ;
    END
  END m_in[86]
  PIN m_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 1096.000 374.350 1100.000 ;
    END
  END m_in[87]
  PIN m_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 1096.000 378.490 1100.000 ;
    END
  END m_in[88]
  PIN m_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 1096.000 382.630 1100.000 ;
    END
  END m_in[89]
  PIN m_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 1096.000 39.930 1100.000 ;
    END
  END m_in[8]
  PIN m_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 1096.000 386.770 1100.000 ;
    END
  END m_in[90]
  PIN m_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 1096.000 391.370 1100.000 ;
    END
  END m_in[91]
  PIN m_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 1096.000 395.510 1100.000 ;
    END
  END m_in[92]
  PIN m_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1096.000 399.650 1100.000 ;
    END
  END m_in[93]
  PIN m_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 1096.000 403.790 1100.000 ;
    END
  END m_in[94]
  PIN m_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 1096.000 407.930 1100.000 ;
    END
  END m_in[95]
  PIN m_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 1096.000 412.530 1100.000 ;
    END
  END m_in[96]
  PIN m_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 1096.000 416.670 1100.000 ;
    END
  END m_in[97]
  PIN m_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 1096.000 420.810 1100.000 ;
    END
  END m_in[98]
  PIN m_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 1096.000 424.950 1100.000 ;
    END
  END m_in[99]
  PIN m_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 1096.000 44.070 1100.000 ;
    END
  END m_in[9]
  PIN m_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 4.120 1100.000 4.720 ;
    END
  END m_out[0]
  PIN m_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 850.040 1100.000 850.640 ;
    END
  END m_out[100]
  PIN m_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 858.880 1100.000 859.480 ;
    END
  END m_out[101]
  PIN m_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 867.040 1100.000 867.640 ;
    END
  END m_out[102]
  PIN m_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 875.200 1100.000 875.800 ;
    END
  END m_out[103]
  PIN m_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 884.040 1100.000 884.640 ;
    END
  END m_out[104]
  PIN m_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 892.200 1100.000 892.800 ;
    END
  END m_out[105]
  PIN m_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 901.040 1100.000 901.640 ;
    END
  END m_out[106]
  PIN m_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 909.200 1100.000 909.800 ;
    END
  END m_out[107]
  PIN m_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 918.040 1100.000 918.640 ;
    END
  END m_out[108]
  PIN m_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 926.200 1100.000 926.800 ;
    END
  END m_out[109]
  PIN m_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 88.440 1100.000 89.040 ;
    END
  END m_out[10]
  PIN m_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 935.040 1100.000 935.640 ;
    END
  END m_out[110]
  PIN m_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 943.200 1100.000 943.800 ;
    END
  END m_out[111]
  PIN m_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 951.360 1100.000 951.960 ;
    END
  END m_out[112]
  PIN m_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 960.200 1100.000 960.800 ;
    END
  END m_out[113]
  PIN m_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 968.360 1100.000 968.960 ;
    END
  END m_out[114]
  PIN m_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 977.200 1100.000 977.800 ;
    END
  END m_out[115]
  PIN m_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 985.360 1100.000 985.960 ;
    END
  END m_out[116]
  PIN m_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 994.200 1100.000 994.800 ;
    END
  END m_out[117]
  PIN m_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1002.360 1100.000 1002.960 ;
    END
  END m_out[118]
  PIN m_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1011.200 1100.000 1011.800 ;
    END
  END m_out[119]
  PIN m_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 96.600 1100.000 97.200 ;
    END
  END m_out[11]
  PIN m_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1019.360 1100.000 1019.960 ;
    END
  END m_out[120]
  PIN m_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1027.520 1100.000 1028.120 ;
    END
  END m_out[121]
  PIN m_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1036.360 1100.000 1036.960 ;
    END
  END m_out[122]
  PIN m_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1044.520 1100.000 1045.120 ;
    END
  END m_out[123]
  PIN m_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1053.360 1100.000 1053.960 ;
    END
  END m_out[124]
  PIN m_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1061.520 1100.000 1062.120 ;
    END
  END m_out[125]
  PIN m_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1070.360 1100.000 1070.960 ;
    END
  END m_out[126]
  PIN m_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1078.520 1100.000 1079.120 ;
    END
  END m_out[127]
  PIN m_out[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1087.360 1100.000 1087.960 ;
    END
  END m_out[128]
  PIN m_out[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1095.520 1100.000 1096.120 ;
    END
  END m_out[129]
  PIN m_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 105.440 1100.000 106.040 ;
    END
  END m_out[12]
  PIN m_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 113.600 1100.000 114.200 ;
    END
  END m_out[13]
  PIN m_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 122.440 1100.000 123.040 ;
    END
  END m_out[14]
  PIN m_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 130.600 1100.000 131.200 ;
    END
  END m_out[15]
  PIN m_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 139.440 1100.000 140.040 ;
    END
  END m_out[16]
  PIN m_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 147.600 1100.000 148.200 ;
    END
  END m_out[17]
  PIN m_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 156.440 1100.000 157.040 ;
    END
  END m_out[18]
  PIN m_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 164.600 1100.000 165.200 ;
    END
  END m_out[19]
  PIN m_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 12.280 1100.000 12.880 ;
    END
  END m_out[1]
  PIN m_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 172.760 1100.000 173.360 ;
    END
  END m_out[20]
  PIN m_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 181.600 1100.000 182.200 ;
    END
  END m_out[21]
  PIN m_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 189.760 1100.000 190.360 ;
    END
  END m_out[22]
  PIN m_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 198.600 1100.000 199.200 ;
    END
  END m_out[23]
  PIN m_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 206.760 1100.000 207.360 ;
    END
  END m_out[24]
  PIN m_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 215.600 1100.000 216.200 ;
    END
  END m_out[25]
  PIN m_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 223.760 1100.000 224.360 ;
    END
  END m_out[26]
  PIN m_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 232.600 1100.000 233.200 ;
    END
  END m_out[27]
  PIN m_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 240.760 1100.000 241.360 ;
    END
  END m_out[28]
  PIN m_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 248.920 1100.000 249.520 ;
    END
  END m_out[29]
  PIN m_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 20.440 1100.000 21.040 ;
    END
  END m_out[2]
  PIN m_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 257.760 1100.000 258.360 ;
    END
  END m_out[30]
  PIN m_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 265.920 1100.000 266.520 ;
    END
  END m_out[31]
  PIN m_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 274.760 1100.000 275.360 ;
    END
  END m_out[32]
  PIN m_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 282.920 1100.000 283.520 ;
    END
  END m_out[33]
  PIN m_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 291.760 1100.000 292.360 ;
    END
  END m_out[34]
  PIN m_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 299.920 1100.000 300.520 ;
    END
  END m_out[35]
  PIN m_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 308.760 1100.000 309.360 ;
    END
  END m_out[36]
  PIN m_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 316.920 1100.000 317.520 ;
    END
  END m_out[37]
  PIN m_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 325.080 1100.000 325.680 ;
    END
  END m_out[38]
  PIN m_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 333.920 1100.000 334.520 ;
    END
  END m_out[39]
  PIN m_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 29.280 1100.000 29.880 ;
    END
  END m_out[3]
  PIN m_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 342.080 1100.000 342.680 ;
    END
  END m_out[40]
  PIN m_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 350.920 1100.000 351.520 ;
    END
  END m_out[41]
  PIN m_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 359.080 1100.000 359.680 ;
    END
  END m_out[42]
  PIN m_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 367.920 1100.000 368.520 ;
    END
  END m_out[43]
  PIN m_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 376.080 1100.000 376.680 ;
    END
  END m_out[44]
  PIN m_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 384.920 1100.000 385.520 ;
    END
  END m_out[45]
  PIN m_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 393.080 1100.000 393.680 ;
    END
  END m_out[46]
  PIN m_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 401.240 1100.000 401.840 ;
    END
  END m_out[47]
  PIN m_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 410.080 1100.000 410.680 ;
    END
  END m_out[48]
  PIN m_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 418.240 1100.000 418.840 ;
    END
  END m_out[49]
  PIN m_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 37.440 1100.000 38.040 ;
    END
  END m_out[4]
  PIN m_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 427.080 1100.000 427.680 ;
    END
  END m_out[50]
  PIN m_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 435.240 1100.000 435.840 ;
    END
  END m_out[51]
  PIN m_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 444.080 1100.000 444.680 ;
    END
  END m_out[52]
  PIN m_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 452.240 1100.000 452.840 ;
    END
  END m_out[53]
  PIN m_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 461.080 1100.000 461.680 ;
    END
  END m_out[54]
  PIN m_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 469.240 1100.000 469.840 ;
    END
  END m_out[55]
  PIN m_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 477.400 1100.000 478.000 ;
    END
  END m_out[56]
  PIN m_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 486.240 1100.000 486.840 ;
    END
  END m_out[57]
  PIN m_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 494.400 1100.000 495.000 ;
    END
  END m_out[58]
  PIN m_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 503.240 1100.000 503.840 ;
    END
  END m_out[59]
  PIN m_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 46.280 1100.000 46.880 ;
    END
  END m_out[5]
  PIN m_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 511.400 1100.000 512.000 ;
    END
  END m_out[60]
  PIN m_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 520.240 1100.000 520.840 ;
    END
  END m_out[61]
  PIN m_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 528.400 1100.000 529.000 ;
    END
  END m_out[62]
  PIN m_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 537.240 1100.000 537.840 ;
    END
  END m_out[63]
  PIN m_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 545.400 1100.000 546.000 ;
    END
  END m_out[64]
  PIN m_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 554.240 1100.000 554.840 ;
    END
  END m_out[65]
  PIN m_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 562.400 1100.000 563.000 ;
    END
  END m_out[66]
  PIN m_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 570.560 1100.000 571.160 ;
    END
  END m_out[67]
  PIN m_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 579.400 1100.000 580.000 ;
    END
  END m_out[68]
  PIN m_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 587.560 1100.000 588.160 ;
    END
  END m_out[69]
  PIN m_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 54.440 1100.000 55.040 ;
    END
  END m_out[6]
  PIN m_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 596.400 1100.000 597.000 ;
    END
  END m_out[70]
  PIN m_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 604.560 1100.000 605.160 ;
    END
  END m_out[71]
  PIN m_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 613.400 1100.000 614.000 ;
    END
  END m_out[72]
  PIN m_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 621.560 1100.000 622.160 ;
    END
  END m_out[73]
  PIN m_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 630.400 1100.000 631.000 ;
    END
  END m_out[74]
  PIN m_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 638.560 1100.000 639.160 ;
    END
  END m_out[75]
  PIN m_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 646.720 1100.000 647.320 ;
    END
  END m_out[76]
  PIN m_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 655.560 1100.000 656.160 ;
    END
  END m_out[77]
  PIN m_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 663.720 1100.000 664.320 ;
    END
  END m_out[78]
  PIN m_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 672.560 1100.000 673.160 ;
    END
  END m_out[79]
  PIN m_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 63.280 1100.000 63.880 ;
    END
  END m_out[7]
  PIN m_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 680.720 1100.000 681.320 ;
    END
  END m_out[80]
  PIN m_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 689.560 1100.000 690.160 ;
    END
  END m_out[81]
  PIN m_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 697.720 1100.000 698.320 ;
    END
  END m_out[82]
  PIN m_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 706.560 1100.000 707.160 ;
    END
  END m_out[83]
  PIN m_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 714.720 1100.000 715.320 ;
    END
  END m_out[84]
  PIN m_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 722.880 1100.000 723.480 ;
    END
  END m_out[85]
  PIN m_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 731.720 1100.000 732.320 ;
    END
  END m_out[86]
  PIN m_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 739.880 1100.000 740.480 ;
    END
  END m_out[87]
  PIN m_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 748.720 1100.000 749.320 ;
    END
  END m_out[88]
  PIN m_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 756.880 1100.000 757.480 ;
    END
  END m_out[89]
  PIN m_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 71.440 1100.000 72.040 ;
    END
  END m_out[8]
  PIN m_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 765.720 1100.000 766.320 ;
    END
  END m_out[90]
  PIN m_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 773.880 1100.000 774.480 ;
    END
  END m_out[91]
  PIN m_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 782.720 1100.000 783.320 ;
    END
  END m_out[92]
  PIN m_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 790.880 1100.000 791.480 ;
    END
  END m_out[93]
  PIN m_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 799.040 1100.000 799.640 ;
    END
  END m_out[94]
  PIN m_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 807.880 1100.000 808.480 ;
    END
  END m_out[95]
  PIN m_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 816.040 1100.000 816.640 ;
    END
  END m_out[96]
  PIN m_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 824.880 1100.000 825.480 ;
    END
  END m_out[97]
  PIN m_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 833.040 1100.000 833.640 ;
    END
  END m_out[98]
  PIN m_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 841.880 1100.000 842.480 ;
    END
  END m_out[99]
  PIN m_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 80.280 1100.000 80.880 ;
    END
  END m_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1094.340 1088.085 ;
      LAYER met1 ;
        RECT 5.520 10.640 1097.490 1098.160 ;
      LAYER met2 ;
        RECT 0.090 1095.720 1.650 1098.190 ;
        RECT 2.490 1095.720 5.790 1098.190 ;
        RECT 6.630 1095.720 9.930 1098.190 ;
        RECT 10.770 1095.720 14.070 1098.190 ;
        RECT 14.910 1095.720 18.210 1098.190 ;
        RECT 19.050 1095.720 22.350 1098.190 ;
        RECT 23.190 1095.720 26.950 1098.190 ;
        RECT 27.790 1095.720 31.090 1098.190 ;
        RECT 31.930 1095.720 35.230 1098.190 ;
        RECT 36.070 1095.720 39.370 1098.190 ;
        RECT 40.210 1095.720 43.510 1098.190 ;
        RECT 44.350 1095.720 48.110 1098.190 ;
        RECT 48.950 1095.720 52.250 1098.190 ;
        RECT 53.090 1095.720 56.390 1098.190 ;
        RECT 57.230 1095.720 60.530 1098.190 ;
        RECT 61.370 1095.720 64.670 1098.190 ;
        RECT 65.510 1095.720 69.270 1098.190 ;
        RECT 70.110 1095.720 73.410 1098.190 ;
        RECT 74.250 1095.720 77.550 1098.190 ;
        RECT 78.390 1095.720 81.690 1098.190 ;
        RECT 82.530 1095.720 85.830 1098.190 ;
        RECT 86.670 1095.720 90.430 1098.190 ;
        RECT 91.270 1095.720 94.570 1098.190 ;
        RECT 95.410 1095.720 98.710 1098.190 ;
        RECT 99.550 1095.720 102.850 1098.190 ;
        RECT 103.690 1095.720 106.990 1098.190 ;
        RECT 107.830 1095.720 111.590 1098.190 ;
        RECT 112.430 1095.720 115.730 1098.190 ;
        RECT 116.570 1095.720 119.870 1098.190 ;
        RECT 120.710 1095.720 124.010 1098.190 ;
        RECT 124.850 1095.720 128.150 1098.190 ;
        RECT 128.990 1095.720 132.750 1098.190 ;
        RECT 133.590 1095.720 136.890 1098.190 ;
        RECT 137.730 1095.720 141.030 1098.190 ;
        RECT 141.870 1095.720 145.170 1098.190 ;
        RECT 146.010 1095.720 149.310 1098.190 ;
        RECT 150.150 1095.720 153.910 1098.190 ;
        RECT 154.750 1095.720 158.050 1098.190 ;
        RECT 158.890 1095.720 162.190 1098.190 ;
        RECT 163.030 1095.720 166.330 1098.190 ;
        RECT 167.170 1095.720 170.470 1098.190 ;
        RECT 171.310 1095.720 175.070 1098.190 ;
        RECT 175.910 1095.720 179.210 1098.190 ;
        RECT 180.050 1095.720 183.350 1098.190 ;
        RECT 184.190 1095.720 187.490 1098.190 ;
        RECT 188.330 1095.720 191.630 1098.190 ;
        RECT 192.470 1095.720 196.230 1098.190 ;
        RECT 197.070 1095.720 200.370 1098.190 ;
        RECT 201.210 1095.720 204.510 1098.190 ;
        RECT 205.350 1095.720 208.650 1098.190 ;
        RECT 209.490 1095.720 212.790 1098.190 ;
        RECT 213.630 1095.720 217.390 1098.190 ;
        RECT 218.230 1095.720 221.530 1098.190 ;
        RECT 222.370 1095.720 225.670 1098.190 ;
        RECT 226.510 1095.720 229.810 1098.190 ;
        RECT 230.650 1095.720 233.950 1098.190 ;
        RECT 234.790 1095.720 238.090 1098.190 ;
        RECT 238.930 1095.720 242.690 1098.190 ;
        RECT 243.530 1095.720 246.830 1098.190 ;
        RECT 247.670 1095.720 250.970 1098.190 ;
        RECT 251.810 1095.720 255.110 1098.190 ;
        RECT 255.950 1095.720 259.250 1098.190 ;
        RECT 260.090 1095.720 263.850 1098.190 ;
        RECT 264.690 1095.720 267.990 1098.190 ;
        RECT 268.830 1095.720 272.130 1098.190 ;
        RECT 272.970 1095.720 276.270 1098.190 ;
        RECT 277.110 1095.720 280.410 1098.190 ;
        RECT 281.250 1095.720 285.010 1098.190 ;
        RECT 285.850 1095.720 289.150 1098.190 ;
        RECT 289.990 1095.720 293.290 1098.190 ;
        RECT 294.130 1095.720 297.430 1098.190 ;
        RECT 298.270 1095.720 301.570 1098.190 ;
        RECT 302.410 1095.720 306.170 1098.190 ;
        RECT 307.010 1095.720 310.310 1098.190 ;
        RECT 311.150 1095.720 314.450 1098.190 ;
        RECT 315.290 1095.720 318.590 1098.190 ;
        RECT 319.430 1095.720 322.730 1098.190 ;
        RECT 323.570 1095.720 327.330 1098.190 ;
        RECT 328.170 1095.720 331.470 1098.190 ;
        RECT 332.310 1095.720 335.610 1098.190 ;
        RECT 336.450 1095.720 339.750 1098.190 ;
        RECT 340.590 1095.720 343.890 1098.190 ;
        RECT 344.730 1095.720 348.490 1098.190 ;
        RECT 349.330 1095.720 352.630 1098.190 ;
        RECT 353.470 1095.720 356.770 1098.190 ;
        RECT 357.610 1095.720 360.910 1098.190 ;
        RECT 361.750 1095.720 365.050 1098.190 ;
        RECT 365.890 1095.720 369.650 1098.190 ;
        RECT 370.490 1095.720 373.790 1098.190 ;
        RECT 374.630 1095.720 377.930 1098.190 ;
        RECT 378.770 1095.720 382.070 1098.190 ;
        RECT 382.910 1095.720 386.210 1098.190 ;
        RECT 387.050 1095.720 390.810 1098.190 ;
        RECT 391.650 1095.720 394.950 1098.190 ;
        RECT 395.790 1095.720 399.090 1098.190 ;
        RECT 399.930 1095.720 403.230 1098.190 ;
        RECT 404.070 1095.720 407.370 1098.190 ;
        RECT 408.210 1095.720 411.970 1098.190 ;
        RECT 412.810 1095.720 416.110 1098.190 ;
        RECT 416.950 1095.720 420.250 1098.190 ;
        RECT 421.090 1095.720 424.390 1098.190 ;
        RECT 425.230 1095.720 428.530 1098.190 ;
        RECT 429.370 1095.720 433.130 1098.190 ;
        RECT 433.970 1095.720 437.270 1098.190 ;
        RECT 438.110 1095.720 441.410 1098.190 ;
        RECT 442.250 1095.720 445.550 1098.190 ;
        RECT 446.390 1095.720 449.690 1098.190 ;
        RECT 450.530 1095.720 453.830 1098.190 ;
        RECT 454.670 1095.720 458.430 1098.190 ;
        RECT 459.270 1095.720 462.570 1098.190 ;
        RECT 463.410 1095.720 466.710 1098.190 ;
        RECT 467.550 1095.720 470.850 1098.190 ;
        RECT 471.690 1095.720 474.990 1098.190 ;
        RECT 475.830 1095.720 479.590 1098.190 ;
        RECT 480.430 1095.720 483.730 1098.190 ;
        RECT 484.570 1095.720 487.870 1098.190 ;
        RECT 488.710 1095.720 492.010 1098.190 ;
        RECT 492.850 1095.720 496.150 1098.190 ;
        RECT 496.990 1095.720 500.750 1098.190 ;
        RECT 501.590 1095.720 504.890 1098.190 ;
        RECT 505.730 1095.720 509.030 1098.190 ;
        RECT 509.870 1095.720 513.170 1098.190 ;
        RECT 514.010 1095.720 517.310 1098.190 ;
        RECT 518.150 1095.720 521.910 1098.190 ;
        RECT 522.750 1095.720 526.050 1098.190 ;
        RECT 526.890 1095.720 530.190 1098.190 ;
        RECT 531.030 1095.720 534.330 1098.190 ;
        RECT 535.170 1095.720 538.470 1098.190 ;
        RECT 539.310 1095.720 543.070 1098.190 ;
        RECT 543.910 1095.720 547.210 1098.190 ;
        RECT 548.050 1095.720 551.350 1098.190 ;
        RECT 552.190 1095.720 555.490 1098.190 ;
        RECT 556.330 1095.720 559.630 1098.190 ;
        RECT 560.470 1095.720 564.230 1098.190 ;
        RECT 565.070 1095.720 568.370 1098.190 ;
        RECT 569.210 1095.720 572.510 1098.190 ;
        RECT 573.350 1095.720 576.650 1098.190 ;
        RECT 577.490 1095.720 580.790 1098.190 ;
        RECT 581.630 1095.720 585.390 1098.190 ;
        RECT 586.230 1095.720 589.530 1098.190 ;
        RECT 590.370 1095.720 593.670 1098.190 ;
        RECT 594.510 1095.720 597.810 1098.190 ;
        RECT 598.650 1095.720 601.950 1098.190 ;
        RECT 602.790 1095.720 606.550 1098.190 ;
        RECT 607.390 1095.720 610.690 1098.190 ;
        RECT 611.530 1095.720 614.830 1098.190 ;
        RECT 615.670 1095.720 618.970 1098.190 ;
        RECT 619.810 1095.720 623.110 1098.190 ;
        RECT 623.950 1095.720 627.710 1098.190 ;
        RECT 628.550 1095.720 631.850 1098.190 ;
        RECT 632.690 1095.720 635.990 1098.190 ;
        RECT 636.830 1095.720 640.130 1098.190 ;
        RECT 640.970 1095.720 644.270 1098.190 ;
        RECT 645.110 1095.720 648.870 1098.190 ;
        RECT 649.710 1095.720 653.010 1098.190 ;
        RECT 653.850 1095.720 657.150 1098.190 ;
        RECT 657.990 1095.720 661.290 1098.190 ;
        RECT 662.130 1095.720 665.430 1098.190 ;
        RECT 666.270 1095.720 669.570 1098.190 ;
        RECT 670.410 1095.720 674.170 1098.190 ;
        RECT 675.010 1095.720 678.310 1098.190 ;
        RECT 679.150 1095.720 682.450 1098.190 ;
        RECT 683.290 1095.720 686.590 1098.190 ;
        RECT 687.430 1095.720 690.730 1098.190 ;
        RECT 691.570 1095.720 695.330 1098.190 ;
        RECT 696.170 1095.720 699.470 1098.190 ;
        RECT 700.310 1095.720 703.610 1098.190 ;
        RECT 704.450 1095.720 707.750 1098.190 ;
        RECT 708.590 1095.720 711.890 1098.190 ;
        RECT 712.730 1095.720 716.490 1098.190 ;
        RECT 717.330 1095.720 720.630 1098.190 ;
        RECT 721.470 1095.720 724.770 1098.190 ;
        RECT 725.610 1095.720 728.910 1098.190 ;
        RECT 729.750 1095.720 733.050 1098.190 ;
        RECT 733.890 1095.720 737.650 1098.190 ;
        RECT 738.490 1095.720 741.790 1098.190 ;
        RECT 742.630 1095.720 745.930 1098.190 ;
        RECT 746.770 1095.720 750.070 1098.190 ;
        RECT 750.910 1095.720 754.210 1098.190 ;
        RECT 755.050 1095.720 758.810 1098.190 ;
        RECT 759.650 1095.720 762.950 1098.190 ;
        RECT 763.790 1095.720 767.090 1098.190 ;
        RECT 767.930 1095.720 771.230 1098.190 ;
        RECT 772.070 1095.720 775.370 1098.190 ;
        RECT 776.210 1095.720 779.970 1098.190 ;
        RECT 780.810 1095.720 784.110 1098.190 ;
        RECT 784.950 1095.720 788.250 1098.190 ;
        RECT 789.090 1095.720 792.390 1098.190 ;
        RECT 793.230 1095.720 796.530 1098.190 ;
        RECT 797.370 1095.720 801.130 1098.190 ;
        RECT 801.970 1095.720 805.270 1098.190 ;
        RECT 806.110 1095.720 809.410 1098.190 ;
        RECT 810.250 1095.720 813.550 1098.190 ;
        RECT 814.390 1095.720 817.690 1098.190 ;
        RECT 818.530 1095.720 822.290 1098.190 ;
        RECT 823.130 1095.720 826.430 1098.190 ;
        RECT 827.270 1095.720 830.570 1098.190 ;
        RECT 831.410 1095.720 834.710 1098.190 ;
        RECT 835.550 1095.720 838.850 1098.190 ;
        RECT 839.690 1095.720 843.450 1098.190 ;
        RECT 844.290 1095.720 847.590 1098.190 ;
        RECT 848.430 1095.720 851.730 1098.190 ;
        RECT 852.570 1095.720 855.870 1098.190 ;
        RECT 856.710 1095.720 860.010 1098.190 ;
        RECT 860.850 1095.720 864.610 1098.190 ;
        RECT 865.450 1095.720 868.750 1098.190 ;
        RECT 869.590 1095.720 872.890 1098.190 ;
        RECT 873.730 1095.720 877.030 1098.190 ;
        RECT 877.870 1095.720 881.170 1098.190 ;
        RECT 882.010 1095.720 885.310 1098.190 ;
        RECT 886.150 1095.720 889.910 1098.190 ;
        RECT 890.750 1095.720 894.050 1098.190 ;
        RECT 894.890 1095.720 898.190 1098.190 ;
        RECT 899.030 1095.720 902.330 1098.190 ;
        RECT 903.170 1095.720 906.470 1098.190 ;
        RECT 907.310 1095.720 911.070 1098.190 ;
        RECT 911.910 1095.720 915.210 1098.190 ;
        RECT 916.050 1095.720 919.350 1098.190 ;
        RECT 920.190 1095.720 923.490 1098.190 ;
        RECT 924.330 1095.720 927.630 1098.190 ;
        RECT 928.470 1095.720 932.230 1098.190 ;
        RECT 933.070 1095.720 936.370 1098.190 ;
        RECT 937.210 1095.720 940.510 1098.190 ;
        RECT 941.350 1095.720 944.650 1098.190 ;
        RECT 945.490 1095.720 948.790 1098.190 ;
        RECT 949.630 1095.720 953.390 1098.190 ;
        RECT 954.230 1095.720 957.530 1098.190 ;
        RECT 958.370 1095.720 961.670 1098.190 ;
        RECT 962.510 1095.720 965.810 1098.190 ;
        RECT 966.650 1095.720 969.950 1098.190 ;
        RECT 970.790 1095.720 974.550 1098.190 ;
        RECT 975.390 1095.720 978.690 1098.190 ;
        RECT 979.530 1095.720 982.830 1098.190 ;
        RECT 983.670 1095.720 986.970 1098.190 ;
        RECT 987.810 1095.720 991.110 1098.190 ;
        RECT 991.950 1095.720 995.710 1098.190 ;
        RECT 996.550 1095.720 999.850 1098.190 ;
        RECT 1000.690 1095.720 1003.990 1098.190 ;
        RECT 1004.830 1095.720 1008.130 1098.190 ;
        RECT 1008.970 1095.720 1012.270 1098.190 ;
        RECT 1013.110 1095.720 1016.870 1098.190 ;
        RECT 1017.710 1095.720 1021.010 1098.190 ;
        RECT 1021.850 1095.720 1025.150 1098.190 ;
        RECT 1025.990 1095.720 1029.290 1098.190 ;
        RECT 1030.130 1095.720 1033.430 1098.190 ;
        RECT 1034.270 1095.720 1038.030 1098.190 ;
        RECT 1038.870 1095.720 1042.170 1098.190 ;
        RECT 1043.010 1095.720 1046.310 1098.190 ;
        RECT 1047.150 1095.720 1050.450 1098.190 ;
        RECT 1051.290 1095.720 1054.590 1098.190 ;
        RECT 1055.430 1095.720 1059.190 1098.190 ;
        RECT 1060.030 1095.720 1063.330 1098.190 ;
        RECT 1064.170 1095.720 1067.470 1098.190 ;
        RECT 1068.310 1095.720 1071.610 1098.190 ;
        RECT 1072.450 1095.720 1075.750 1098.190 ;
        RECT 1076.590 1095.720 1080.350 1098.190 ;
        RECT 1081.190 1095.720 1084.490 1098.190 ;
        RECT 1085.330 1095.720 1088.630 1098.190 ;
        RECT 1089.470 1095.720 1092.770 1098.190 ;
        RECT 1093.610 1095.720 1096.910 1098.190 ;
        RECT 0.090 4.235 1097.460 1095.720 ;
      LAYER met3 ;
        RECT 0.065 1095.120 1095.600 1095.985 ;
        RECT 0.065 1088.360 1096.000 1095.120 ;
        RECT 0.065 1086.960 1095.600 1088.360 ;
        RECT 0.065 1079.520 1096.000 1086.960 ;
        RECT 0.065 1078.120 1095.600 1079.520 ;
        RECT 0.065 1071.360 1096.000 1078.120 ;
        RECT 0.065 1069.960 1095.600 1071.360 ;
        RECT 0.065 1062.520 1096.000 1069.960 ;
        RECT 0.065 1061.120 1095.600 1062.520 ;
        RECT 0.065 1054.360 1096.000 1061.120 ;
        RECT 0.065 1052.960 1095.600 1054.360 ;
        RECT 0.065 1045.520 1096.000 1052.960 ;
        RECT 0.065 1044.120 1095.600 1045.520 ;
        RECT 0.065 1037.360 1096.000 1044.120 ;
        RECT 0.065 1035.960 1095.600 1037.360 ;
        RECT 0.065 1028.520 1096.000 1035.960 ;
        RECT 0.065 1027.120 1095.600 1028.520 ;
        RECT 0.065 1020.360 1096.000 1027.120 ;
        RECT 0.065 1018.960 1095.600 1020.360 ;
        RECT 0.065 1012.200 1096.000 1018.960 ;
        RECT 0.065 1010.800 1095.600 1012.200 ;
        RECT 0.065 1003.360 1096.000 1010.800 ;
        RECT 0.065 1001.960 1095.600 1003.360 ;
        RECT 0.065 995.200 1096.000 1001.960 ;
        RECT 0.065 993.800 1095.600 995.200 ;
        RECT 0.065 986.360 1096.000 993.800 ;
        RECT 0.065 984.960 1095.600 986.360 ;
        RECT 0.065 978.200 1096.000 984.960 ;
        RECT 0.065 976.800 1095.600 978.200 ;
        RECT 0.065 969.360 1096.000 976.800 ;
        RECT 0.065 967.960 1095.600 969.360 ;
        RECT 0.065 961.200 1096.000 967.960 ;
        RECT 0.065 959.800 1095.600 961.200 ;
        RECT 0.065 952.360 1096.000 959.800 ;
        RECT 0.065 950.960 1095.600 952.360 ;
        RECT 0.065 944.200 1096.000 950.960 ;
        RECT 0.065 942.800 1095.600 944.200 ;
        RECT 0.065 936.040 1096.000 942.800 ;
        RECT 0.065 934.640 1095.600 936.040 ;
        RECT 0.065 927.200 1096.000 934.640 ;
        RECT 0.065 925.800 1095.600 927.200 ;
        RECT 0.065 919.040 1096.000 925.800 ;
        RECT 0.065 917.640 1095.600 919.040 ;
        RECT 0.065 910.200 1096.000 917.640 ;
        RECT 0.065 908.800 1095.600 910.200 ;
        RECT 0.065 902.040 1096.000 908.800 ;
        RECT 0.065 900.640 1095.600 902.040 ;
        RECT 0.065 893.200 1096.000 900.640 ;
        RECT 0.065 891.800 1095.600 893.200 ;
        RECT 0.065 885.040 1096.000 891.800 ;
        RECT 0.065 883.640 1095.600 885.040 ;
        RECT 0.065 876.200 1096.000 883.640 ;
        RECT 0.065 874.800 1095.600 876.200 ;
        RECT 0.065 868.040 1096.000 874.800 ;
        RECT 0.065 866.640 1095.600 868.040 ;
        RECT 0.065 859.880 1096.000 866.640 ;
        RECT 0.065 858.480 1095.600 859.880 ;
        RECT 0.065 851.040 1096.000 858.480 ;
        RECT 0.065 849.640 1095.600 851.040 ;
        RECT 0.065 842.880 1096.000 849.640 ;
        RECT 0.065 841.480 1095.600 842.880 ;
        RECT 0.065 834.040 1096.000 841.480 ;
        RECT 0.065 832.640 1095.600 834.040 ;
        RECT 0.065 825.880 1096.000 832.640 ;
        RECT 0.065 824.480 1095.600 825.880 ;
        RECT 0.065 817.040 1096.000 824.480 ;
        RECT 0.065 815.640 1095.600 817.040 ;
        RECT 0.065 808.880 1096.000 815.640 ;
        RECT 0.065 807.480 1095.600 808.880 ;
        RECT 0.065 800.040 1096.000 807.480 ;
        RECT 0.065 798.640 1095.600 800.040 ;
        RECT 0.065 791.880 1096.000 798.640 ;
        RECT 0.065 790.480 1095.600 791.880 ;
        RECT 0.065 783.720 1096.000 790.480 ;
        RECT 0.065 782.320 1095.600 783.720 ;
        RECT 0.065 774.880 1096.000 782.320 ;
        RECT 0.065 773.480 1095.600 774.880 ;
        RECT 0.065 766.720 1096.000 773.480 ;
        RECT 0.065 765.320 1095.600 766.720 ;
        RECT 0.065 757.880 1096.000 765.320 ;
        RECT 0.065 756.480 1095.600 757.880 ;
        RECT 0.065 749.720 1096.000 756.480 ;
        RECT 0.065 748.320 1095.600 749.720 ;
        RECT 0.065 740.880 1096.000 748.320 ;
        RECT 0.065 739.480 1095.600 740.880 ;
        RECT 0.065 732.720 1096.000 739.480 ;
        RECT 0.065 731.320 1095.600 732.720 ;
        RECT 0.065 723.880 1096.000 731.320 ;
        RECT 0.065 722.480 1095.600 723.880 ;
        RECT 0.065 715.720 1096.000 722.480 ;
        RECT 0.065 714.320 1095.600 715.720 ;
        RECT 0.065 707.560 1096.000 714.320 ;
        RECT 0.065 706.160 1095.600 707.560 ;
        RECT 0.065 698.720 1096.000 706.160 ;
        RECT 0.065 697.320 1095.600 698.720 ;
        RECT 0.065 690.560 1096.000 697.320 ;
        RECT 0.065 689.160 1095.600 690.560 ;
        RECT 0.065 681.720 1096.000 689.160 ;
        RECT 0.065 680.320 1095.600 681.720 ;
        RECT 0.065 673.560 1096.000 680.320 ;
        RECT 0.065 672.160 1095.600 673.560 ;
        RECT 0.065 664.720 1096.000 672.160 ;
        RECT 0.065 663.320 1095.600 664.720 ;
        RECT 0.065 656.560 1096.000 663.320 ;
        RECT 0.065 655.160 1095.600 656.560 ;
        RECT 0.065 647.720 1096.000 655.160 ;
        RECT 0.065 646.320 1095.600 647.720 ;
        RECT 0.065 639.560 1096.000 646.320 ;
        RECT 0.065 638.160 1095.600 639.560 ;
        RECT 0.065 631.400 1096.000 638.160 ;
        RECT 0.065 630.000 1095.600 631.400 ;
        RECT 0.065 622.560 1096.000 630.000 ;
        RECT 0.065 621.160 1095.600 622.560 ;
        RECT 0.065 614.400 1096.000 621.160 ;
        RECT 0.065 613.000 1095.600 614.400 ;
        RECT 0.065 605.560 1096.000 613.000 ;
        RECT 0.065 604.160 1095.600 605.560 ;
        RECT 0.065 597.400 1096.000 604.160 ;
        RECT 0.065 596.000 1095.600 597.400 ;
        RECT 0.065 588.560 1096.000 596.000 ;
        RECT 0.065 587.160 1095.600 588.560 ;
        RECT 0.065 580.400 1096.000 587.160 ;
        RECT 0.065 579.000 1095.600 580.400 ;
        RECT 0.065 571.560 1096.000 579.000 ;
        RECT 0.065 570.160 1095.600 571.560 ;
        RECT 0.065 563.400 1096.000 570.160 ;
        RECT 0.065 562.000 1095.600 563.400 ;
        RECT 0.065 555.240 1096.000 562.000 ;
        RECT 0.065 553.840 1095.600 555.240 ;
        RECT 0.065 546.400 1096.000 553.840 ;
        RECT 0.065 545.000 1095.600 546.400 ;
        RECT 0.065 538.240 1096.000 545.000 ;
        RECT 0.065 536.840 1095.600 538.240 ;
        RECT 0.065 529.400 1096.000 536.840 ;
        RECT 0.065 528.000 1095.600 529.400 ;
        RECT 0.065 521.240 1096.000 528.000 ;
        RECT 0.065 519.840 1095.600 521.240 ;
        RECT 0.065 512.400 1096.000 519.840 ;
        RECT 0.065 511.000 1095.600 512.400 ;
        RECT 0.065 504.240 1096.000 511.000 ;
        RECT 0.065 502.840 1095.600 504.240 ;
        RECT 0.065 495.400 1096.000 502.840 ;
        RECT 0.065 494.000 1095.600 495.400 ;
        RECT 0.065 487.240 1096.000 494.000 ;
        RECT 0.065 485.840 1095.600 487.240 ;
        RECT 0.065 478.400 1096.000 485.840 ;
        RECT 0.065 477.000 1095.600 478.400 ;
        RECT 0.065 470.240 1096.000 477.000 ;
        RECT 0.065 468.840 1095.600 470.240 ;
        RECT 0.065 462.080 1096.000 468.840 ;
        RECT 0.065 460.680 1095.600 462.080 ;
        RECT 0.065 453.240 1096.000 460.680 ;
        RECT 0.065 451.840 1095.600 453.240 ;
        RECT 0.065 445.080 1096.000 451.840 ;
        RECT 0.065 443.680 1095.600 445.080 ;
        RECT 0.065 436.240 1096.000 443.680 ;
        RECT 0.065 434.840 1095.600 436.240 ;
        RECT 0.065 428.080 1096.000 434.840 ;
        RECT 0.065 426.680 1095.600 428.080 ;
        RECT 0.065 419.240 1096.000 426.680 ;
        RECT 0.065 417.840 1095.600 419.240 ;
        RECT 0.065 411.080 1096.000 417.840 ;
        RECT 0.065 409.680 1095.600 411.080 ;
        RECT 0.065 402.240 1096.000 409.680 ;
        RECT 0.065 400.840 1095.600 402.240 ;
        RECT 0.065 394.080 1096.000 400.840 ;
        RECT 0.065 392.680 1095.600 394.080 ;
        RECT 0.065 385.920 1096.000 392.680 ;
        RECT 0.065 384.520 1095.600 385.920 ;
        RECT 0.065 377.080 1096.000 384.520 ;
        RECT 0.065 375.680 1095.600 377.080 ;
        RECT 0.065 368.920 1096.000 375.680 ;
        RECT 0.065 367.520 1095.600 368.920 ;
        RECT 0.065 360.080 1096.000 367.520 ;
        RECT 0.065 358.680 1095.600 360.080 ;
        RECT 0.065 351.920 1096.000 358.680 ;
        RECT 0.065 350.520 1095.600 351.920 ;
        RECT 0.065 343.080 1096.000 350.520 ;
        RECT 0.065 341.680 1095.600 343.080 ;
        RECT 0.065 334.920 1096.000 341.680 ;
        RECT 0.065 333.520 1095.600 334.920 ;
        RECT 0.065 326.080 1096.000 333.520 ;
        RECT 0.065 324.680 1095.600 326.080 ;
        RECT 0.065 317.920 1096.000 324.680 ;
        RECT 0.065 316.520 1095.600 317.920 ;
        RECT 0.065 309.760 1096.000 316.520 ;
        RECT 0.065 308.360 1095.600 309.760 ;
        RECT 0.065 300.920 1096.000 308.360 ;
        RECT 0.065 299.520 1095.600 300.920 ;
        RECT 0.065 292.760 1096.000 299.520 ;
        RECT 0.065 291.360 1095.600 292.760 ;
        RECT 0.065 283.920 1096.000 291.360 ;
        RECT 0.065 282.520 1095.600 283.920 ;
        RECT 0.065 275.760 1096.000 282.520 ;
        RECT 0.065 274.360 1095.600 275.760 ;
        RECT 0.065 266.920 1096.000 274.360 ;
        RECT 0.065 265.520 1095.600 266.920 ;
        RECT 0.065 258.760 1096.000 265.520 ;
        RECT 0.065 257.360 1095.600 258.760 ;
        RECT 0.065 249.920 1096.000 257.360 ;
        RECT 0.065 248.520 1095.600 249.920 ;
        RECT 0.065 241.760 1096.000 248.520 ;
        RECT 0.065 240.360 1095.600 241.760 ;
        RECT 0.065 233.600 1096.000 240.360 ;
        RECT 0.065 232.200 1095.600 233.600 ;
        RECT 0.065 224.760 1096.000 232.200 ;
        RECT 0.065 223.360 1095.600 224.760 ;
        RECT 0.065 216.600 1096.000 223.360 ;
        RECT 0.065 215.200 1095.600 216.600 ;
        RECT 0.065 207.760 1096.000 215.200 ;
        RECT 0.065 206.360 1095.600 207.760 ;
        RECT 0.065 199.600 1096.000 206.360 ;
        RECT 0.065 198.200 1095.600 199.600 ;
        RECT 0.065 190.760 1096.000 198.200 ;
        RECT 0.065 189.360 1095.600 190.760 ;
        RECT 0.065 182.600 1096.000 189.360 ;
        RECT 0.065 181.200 1095.600 182.600 ;
        RECT 0.065 173.760 1096.000 181.200 ;
        RECT 0.065 172.360 1095.600 173.760 ;
        RECT 0.065 165.600 1096.000 172.360 ;
        RECT 0.065 164.200 1095.600 165.600 ;
        RECT 0.065 157.440 1096.000 164.200 ;
        RECT 0.065 156.040 1095.600 157.440 ;
        RECT 0.065 148.600 1096.000 156.040 ;
        RECT 0.065 147.200 1095.600 148.600 ;
        RECT 0.065 140.440 1096.000 147.200 ;
        RECT 0.065 139.040 1095.600 140.440 ;
        RECT 0.065 131.600 1096.000 139.040 ;
        RECT 0.065 130.200 1095.600 131.600 ;
        RECT 0.065 123.440 1096.000 130.200 ;
        RECT 0.065 122.040 1095.600 123.440 ;
        RECT 0.065 114.600 1096.000 122.040 ;
        RECT 0.065 113.200 1095.600 114.600 ;
        RECT 0.065 106.440 1096.000 113.200 ;
        RECT 0.065 105.040 1095.600 106.440 ;
        RECT 0.065 97.600 1096.000 105.040 ;
        RECT 0.065 96.200 1095.600 97.600 ;
        RECT 0.065 89.440 1096.000 96.200 ;
        RECT 0.065 88.040 1095.600 89.440 ;
        RECT 0.065 81.280 1096.000 88.040 ;
        RECT 0.065 79.880 1095.600 81.280 ;
        RECT 0.065 72.440 1096.000 79.880 ;
        RECT 0.065 71.040 1095.600 72.440 ;
        RECT 0.065 64.280 1096.000 71.040 ;
        RECT 0.065 62.880 1095.600 64.280 ;
        RECT 0.065 55.440 1096.000 62.880 ;
        RECT 0.065 54.040 1095.600 55.440 ;
        RECT 0.065 47.280 1096.000 54.040 ;
        RECT 0.065 45.880 1095.600 47.280 ;
        RECT 0.065 38.440 1096.000 45.880 ;
        RECT 0.065 37.040 1095.600 38.440 ;
        RECT 0.065 30.280 1096.000 37.040 ;
        RECT 0.065 28.880 1095.600 30.280 ;
        RECT 0.065 21.440 1096.000 28.880 ;
        RECT 0.065 20.040 1095.600 21.440 ;
        RECT 0.065 13.280 1096.000 20.040 ;
        RECT 0.065 11.880 1095.600 13.280 ;
        RECT 0.065 5.120 1096.000 11.880 ;
        RECT 0.065 4.255 1095.600 5.120 ;
      LAYER met4 ;
        RECT 17.775 68.855 20.640 1085.785 ;
        RECT 23.040 68.855 97.440 1085.785 ;
        RECT 99.840 68.855 174.240 1085.785 ;
        RECT 176.640 68.855 251.040 1085.785 ;
        RECT 253.440 68.855 327.840 1085.785 ;
        RECT 330.240 68.855 404.640 1085.785 ;
        RECT 407.040 68.855 481.440 1085.785 ;
        RECT 483.840 68.855 558.240 1085.785 ;
        RECT 560.640 68.855 635.040 1085.785 ;
        RECT 637.440 68.855 711.840 1085.785 ;
        RECT 714.240 68.855 788.640 1085.785 ;
        RECT 791.040 68.855 865.440 1085.785 ;
        RECT 867.840 68.855 942.240 1085.785 ;
        RECT 944.640 68.855 1019.040 1085.785 ;
        RECT 1021.440 68.855 1089.905 1085.785 ;
  END
END multiply_4
END LIBRARY

