VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO icache
  CLASS BLOCK ;
  FOREIGN icache ;
  ORIGIN 0.000 0.000 ;
  SIZE 680.000 BY 680.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 2.080 680.000 2.680 ;
    END
  END clk
  PIN flush_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END flush_in
  PIN i_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END i_in[0]
  PIN i_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END i_in[10]
  PIN i_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END i_in[11]
  PIN i_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END i_in[12]
  PIN i_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END i_in[13]
  PIN i_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END i_in[14]
  PIN i_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END i_in[15]
  PIN i_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END i_in[16]
  PIN i_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END i_in[17]
  PIN i_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END i_in[18]
  PIN i_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END i_in[19]
  PIN i_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END i_in[1]
  PIN i_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END i_in[20]
  PIN i_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END i_in[21]
  PIN i_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END i_in[22]
  PIN i_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END i_in[23]
  PIN i_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END i_in[24]
  PIN i_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END i_in[25]
  PIN i_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END i_in[26]
  PIN i_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END i_in[27]
  PIN i_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END i_in[28]
  PIN i_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END i_in[29]
  PIN i_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END i_in[2]
  PIN i_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END i_in[30]
  PIN i_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END i_in[31]
  PIN i_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END i_in[32]
  PIN i_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END i_in[33]
  PIN i_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END i_in[34]
  PIN i_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END i_in[35]
  PIN i_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END i_in[36]
  PIN i_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END i_in[37]
  PIN i_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END i_in[38]
  PIN i_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END i_in[39]
  PIN i_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END i_in[3]
  PIN i_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END i_in[40]
  PIN i_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END i_in[41]
  PIN i_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END i_in[42]
  PIN i_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END i_in[43]
  PIN i_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END i_in[44]
  PIN i_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END i_in[45]
  PIN i_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END i_in[46]
  PIN i_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END i_in[47]
  PIN i_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END i_in[48]
  PIN i_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END i_in[49]
  PIN i_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END i_in[4]
  PIN i_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END i_in[50]
  PIN i_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END i_in[51]
  PIN i_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END i_in[52]
  PIN i_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END i_in[53]
  PIN i_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END i_in[54]
  PIN i_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END i_in[55]
  PIN i_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END i_in[56]
  PIN i_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END i_in[57]
  PIN i_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END i_in[58]
  PIN i_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END i_in[59]
  PIN i_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END i_in[5]
  PIN i_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END i_in[60]
  PIN i_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END i_in[61]
  PIN i_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END i_in[62]
  PIN i_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END i_in[63]
  PIN i_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END i_in[64]
  PIN i_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END i_in[65]
  PIN i_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END i_in[66]
  PIN i_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END i_in[67]
  PIN i_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END i_in[68]
  PIN i_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END i_in[69]
  PIN i_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END i_in[6]
  PIN i_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END i_in[7]
  PIN i_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END i_in[8]
  PIN i_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END i_in[9]
  PIN i_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END i_out[0]
  PIN i_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END i_out[10]
  PIN i_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END i_out[11]
  PIN i_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END i_out[12]
  PIN i_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END i_out[13]
  PIN i_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END i_out[14]
  PIN i_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END i_out[15]
  PIN i_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END i_out[16]
  PIN i_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END i_out[17]
  PIN i_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END i_out[18]
  PIN i_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END i_out[19]
  PIN i_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END i_out[1]
  PIN i_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END i_out[20]
  PIN i_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END i_out[21]
  PIN i_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END i_out[22]
  PIN i_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END i_out[23]
  PIN i_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END i_out[24]
  PIN i_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END i_out[25]
  PIN i_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END i_out[26]
  PIN i_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END i_out[27]
  PIN i_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END i_out[28]
  PIN i_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END i_out[29]
  PIN i_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END i_out[2]
  PIN i_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END i_out[30]
  PIN i_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END i_out[31]
  PIN i_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END i_out[32]
  PIN i_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END i_out[33]
  PIN i_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END i_out[34]
  PIN i_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END i_out[35]
  PIN i_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END i_out[36]
  PIN i_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END i_out[37]
  PIN i_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END i_out[38]
  PIN i_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END i_out[39]
  PIN i_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END i_out[3]
  PIN i_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 4.000 ;
    END
  END i_out[40]
  PIN i_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END i_out[41]
  PIN i_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END i_out[42]
  PIN i_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END i_out[43]
  PIN i_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END i_out[44]
  PIN i_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END i_out[45]
  PIN i_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END i_out[46]
  PIN i_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END i_out[47]
  PIN i_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END i_out[48]
  PIN i_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END i_out[49]
  PIN i_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END i_out[4]
  PIN i_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END i_out[50]
  PIN i_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END i_out[51]
  PIN i_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END i_out[52]
  PIN i_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END i_out[53]
  PIN i_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END i_out[54]
  PIN i_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END i_out[55]
  PIN i_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END i_out[56]
  PIN i_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END i_out[57]
  PIN i_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END i_out[58]
  PIN i_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END i_out[59]
  PIN i_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END i_out[5]
  PIN i_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END i_out[60]
  PIN i_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 0.000 516.950 4.000 ;
    END
  END i_out[61]
  PIN i_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END i_out[62]
  PIN i_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END i_out[63]
  PIN i_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END i_out[64]
  PIN i_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END i_out[65]
  PIN i_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END i_out[66]
  PIN i_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END i_out[67]
  PIN i_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END i_out[68]
  PIN i_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END i_out[69]
  PIN i_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END i_out[6]
  PIN i_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END i_out[70]
  PIN i_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END i_out[71]
  PIN i_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END i_out[72]
  PIN i_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END i_out[73]
  PIN i_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END i_out[74]
  PIN i_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END i_out[75]
  PIN i_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END i_out[76]
  PIN i_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END i_out[77]
  PIN i_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END i_out[78]
  PIN i_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END i_out[79]
  PIN i_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END i_out[7]
  PIN i_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END i_out[80]
  PIN i_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END i_out[81]
  PIN i_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END i_out[82]
  PIN i_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END i_out[83]
  PIN i_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END i_out[84]
  PIN i_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END i_out[85]
  PIN i_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END i_out[86]
  PIN i_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END i_out[87]
  PIN i_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END i_out[88]
  PIN i_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END i_out[89]
  PIN i_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END i_out[8]
  PIN i_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END i_out[90]
  PIN i_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END i_out[91]
  PIN i_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END i_out[92]
  PIN i_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 0.000 642.530 4.000 ;
    END
  END i_out[93]
  PIN i_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END i_out[94]
  PIN i_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END i_out[95]
  PIN i_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END i_out[96]
  PIN i_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END i_out[97]
  PIN i_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 0.000 662.310 4.000 ;
    END
  END i_out[98]
  PIN i_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END i_out[9]
  PIN inval_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END inval_in
  PIN m_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 12.280 680.000 12.880 ;
    END
  END m_in[0]
  PIN m_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 522.960 680.000 523.560 ;
    END
  END m_in[100]
  PIN m_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 528.400 680.000 529.000 ;
    END
  END m_in[101]
  PIN m_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 533.160 680.000 533.760 ;
    END
  END m_in[102]
  PIN m_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 538.600 680.000 539.200 ;
    END
  END m_in[103]
  PIN m_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 543.360 680.000 543.960 ;
    END
  END m_in[104]
  PIN m_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 548.800 680.000 549.400 ;
    END
  END m_in[105]
  PIN m_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 554.240 680.000 554.840 ;
    END
  END m_in[106]
  PIN m_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 559.000 680.000 559.600 ;
    END
  END m_in[107]
  PIN m_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 564.440 680.000 565.040 ;
    END
  END m_in[108]
  PIN m_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 569.200 680.000 569.800 ;
    END
  END m_in[109]
  PIN m_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 63.280 680.000 63.880 ;
    END
  END m_in[10]
  PIN m_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 574.640 680.000 575.240 ;
    END
  END m_in[110]
  PIN m_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 579.400 680.000 580.000 ;
    END
  END m_in[111]
  PIN m_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 584.840 680.000 585.440 ;
    END
  END m_in[112]
  PIN m_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 589.600 680.000 590.200 ;
    END
  END m_in[113]
  PIN m_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 595.040 680.000 595.640 ;
    END
  END m_in[114]
  PIN m_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 599.800 680.000 600.400 ;
    END
  END m_in[115]
  PIN m_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 605.240 680.000 605.840 ;
    END
  END m_in[116]
  PIN m_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 610.000 680.000 610.600 ;
    END
  END m_in[117]
  PIN m_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 615.440 680.000 616.040 ;
    END
  END m_in[118]
  PIN m_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 620.200 680.000 620.800 ;
    END
  END m_in[119]
  PIN m_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 68.040 680.000 68.640 ;
    END
  END m_in[11]
  PIN m_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 625.640 680.000 626.240 ;
    END
  END m_in[120]
  PIN m_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 630.400 680.000 631.000 ;
    END
  END m_in[121]
  PIN m_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 635.840 680.000 636.440 ;
    END
  END m_in[122]
  PIN m_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 640.600 680.000 641.200 ;
    END
  END m_in[123]
  PIN m_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 646.040 680.000 646.640 ;
    END
  END m_in[124]
  PIN m_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 650.800 680.000 651.400 ;
    END
  END m_in[125]
  PIN m_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 656.240 680.000 656.840 ;
    END
  END m_in[126]
  PIN m_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 661.000 680.000 661.600 ;
    END
  END m_in[127]
  PIN m_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 666.440 680.000 667.040 ;
    END
  END m_in[128]
  PIN m_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 671.200 680.000 671.800 ;
    END
  END m_in[129]
  PIN m_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 73.480 680.000 74.080 ;
    END
  END m_in[12]
  PIN m_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 676.640 680.000 677.240 ;
    END
  END m_in[130]
  PIN m_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 78.240 680.000 78.840 ;
    END
  END m_in[13]
  PIN m_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 83.680 680.000 84.280 ;
    END
  END m_in[14]
  PIN m_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 88.440 680.000 89.040 ;
    END
  END m_in[15]
  PIN m_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 93.880 680.000 94.480 ;
    END
  END m_in[16]
  PIN m_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 98.640 680.000 99.240 ;
    END
  END m_in[17]
  PIN m_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 104.080 680.000 104.680 ;
    END
  END m_in[18]
  PIN m_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 108.840 680.000 109.440 ;
    END
  END m_in[19]
  PIN m_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 17.040 680.000 17.640 ;
    END
  END m_in[1]
  PIN m_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 114.280 680.000 114.880 ;
    END
  END m_in[20]
  PIN m_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 119.040 680.000 119.640 ;
    END
  END m_in[21]
  PIN m_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 124.480 680.000 125.080 ;
    END
  END m_in[22]
  PIN m_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 129.240 680.000 129.840 ;
    END
  END m_in[23]
  PIN m_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 134.680 680.000 135.280 ;
    END
  END m_in[24]
  PIN m_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 140.120 680.000 140.720 ;
    END
  END m_in[25]
  PIN m_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 144.880 680.000 145.480 ;
    END
  END m_in[26]
  PIN m_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 150.320 680.000 150.920 ;
    END
  END m_in[27]
  PIN m_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 155.080 680.000 155.680 ;
    END
  END m_in[28]
  PIN m_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 160.520 680.000 161.120 ;
    END
  END m_in[29]
  PIN m_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 22.480 680.000 23.080 ;
    END
  END m_in[2]
  PIN m_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 165.280 680.000 165.880 ;
    END
  END m_in[30]
  PIN m_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 170.720 680.000 171.320 ;
    END
  END m_in[31]
  PIN m_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 175.480 680.000 176.080 ;
    END
  END m_in[32]
  PIN m_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 180.920 680.000 181.520 ;
    END
  END m_in[33]
  PIN m_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 185.680 680.000 186.280 ;
    END
  END m_in[34]
  PIN m_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 191.120 680.000 191.720 ;
    END
  END m_in[35]
  PIN m_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 195.880 680.000 196.480 ;
    END
  END m_in[36]
  PIN m_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 201.320 680.000 201.920 ;
    END
  END m_in[37]
  PIN m_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 206.080 680.000 206.680 ;
    END
  END m_in[38]
  PIN m_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 211.520 680.000 212.120 ;
    END
  END m_in[39]
  PIN m_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 27.240 680.000 27.840 ;
    END
  END m_in[3]
  PIN m_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 216.280 680.000 216.880 ;
    END
  END m_in[40]
  PIN m_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 221.720 680.000 222.320 ;
    END
  END m_in[41]
  PIN m_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 226.480 680.000 227.080 ;
    END
  END m_in[42]
  PIN m_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 231.920 680.000 232.520 ;
    END
  END m_in[43]
  PIN m_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 236.680 680.000 237.280 ;
    END
  END m_in[44]
  PIN m_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 242.120 680.000 242.720 ;
    END
  END m_in[45]
  PIN m_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 246.880 680.000 247.480 ;
    END
  END m_in[46]
  PIN m_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 252.320 680.000 252.920 ;
    END
  END m_in[47]
  PIN m_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 257.080 680.000 257.680 ;
    END
  END m_in[48]
  PIN m_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 262.520 680.000 263.120 ;
    END
  END m_in[49]
  PIN m_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 32.680 680.000 33.280 ;
    END
  END m_in[4]
  PIN m_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 267.280 680.000 267.880 ;
    END
  END m_in[50]
  PIN m_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 272.720 680.000 273.320 ;
    END
  END m_in[51]
  PIN m_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 278.160 680.000 278.760 ;
    END
  END m_in[52]
  PIN m_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 282.920 680.000 283.520 ;
    END
  END m_in[53]
  PIN m_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 288.360 680.000 288.960 ;
    END
  END m_in[54]
  PIN m_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 293.120 680.000 293.720 ;
    END
  END m_in[55]
  PIN m_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 298.560 680.000 299.160 ;
    END
  END m_in[56]
  PIN m_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 303.320 680.000 303.920 ;
    END
  END m_in[57]
  PIN m_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 308.760 680.000 309.360 ;
    END
  END m_in[58]
  PIN m_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 313.520 680.000 314.120 ;
    END
  END m_in[59]
  PIN m_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 37.440 680.000 38.040 ;
    END
  END m_in[5]
  PIN m_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 318.960 680.000 319.560 ;
    END
  END m_in[60]
  PIN m_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 323.720 680.000 324.320 ;
    END
  END m_in[61]
  PIN m_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 329.160 680.000 329.760 ;
    END
  END m_in[62]
  PIN m_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 333.920 680.000 334.520 ;
    END
  END m_in[63]
  PIN m_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 339.360 680.000 339.960 ;
    END
  END m_in[64]
  PIN m_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 344.120 680.000 344.720 ;
    END
  END m_in[65]
  PIN m_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 349.560 680.000 350.160 ;
    END
  END m_in[66]
  PIN m_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 354.320 680.000 354.920 ;
    END
  END m_in[67]
  PIN m_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 359.760 680.000 360.360 ;
    END
  END m_in[68]
  PIN m_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 364.520 680.000 365.120 ;
    END
  END m_in[69]
  PIN m_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 42.880 680.000 43.480 ;
    END
  END m_in[6]
  PIN m_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 369.960 680.000 370.560 ;
    END
  END m_in[70]
  PIN m_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 374.720 680.000 375.320 ;
    END
  END m_in[71]
  PIN m_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 380.160 680.000 380.760 ;
    END
  END m_in[72]
  PIN m_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 384.920 680.000 385.520 ;
    END
  END m_in[73]
  PIN m_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 390.360 680.000 390.960 ;
    END
  END m_in[74]
  PIN m_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 395.120 680.000 395.720 ;
    END
  END m_in[75]
  PIN m_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 400.560 680.000 401.160 ;
    END
  END m_in[76]
  PIN m_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 405.320 680.000 405.920 ;
    END
  END m_in[77]
  PIN m_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 410.760 680.000 411.360 ;
    END
  END m_in[78]
  PIN m_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 416.200 680.000 416.800 ;
    END
  END m_in[79]
  PIN m_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 47.640 680.000 48.240 ;
    END
  END m_in[7]
  PIN m_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 420.960 680.000 421.560 ;
    END
  END m_in[80]
  PIN m_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 426.400 680.000 427.000 ;
    END
  END m_in[81]
  PIN m_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 431.160 680.000 431.760 ;
    END
  END m_in[82]
  PIN m_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 436.600 680.000 437.200 ;
    END
  END m_in[83]
  PIN m_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 441.360 680.000 441.960 ;
    END
  END m_in[84]
  PIN m_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 446.800 680.000 447.400 ;
    END
  END m_in[85]
  PIN m_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 451.560 680.000 452.160 ;
    END
  END m_in[86]
  PIN m_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 457.000 680.000 457.600 ;
    END
  END m_in[87]
  PIN m_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 461.760 680.000 462.360 ;
    END
  END m_in[88]
  PIN m_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 467.200 680.000 467.800 ;
    END
  END m_in[89]
  PIN m_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 53.080 680.000 53.680 ;
    END
  END m_in[8]
  PIN m_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 471.960 680.000 472.560 ;
    END
  END m_in[90]
  PIN m_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 477.400 680.000 478.000 ;
    END
  END m_in[91]
  PIN m_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 482.160 680.000 482.760 ;
    END
  END m_in[92]
  PIN m_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 487.600 680.000 488.200 ;
    END
  END m_in[93]
  PIN m_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 492.360 680.000 492.960 ;
    END
  END m_in[94]
  PIN m_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 497.800 680.000 498.400 ;
    END
  END m_in[95]
  PIN m_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 502.560 680.000 503.160 ;
    END
  END m_in[96]
  PIN m_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 508.000 680.000 508.600 ;
    END
  END m_in[97]
  PIN m_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 512.760 680.000 513.360 ;
    END
  END m_in[98]
  PIN m_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 518.200 680.000 518.800 ;
    END
  END m_in[99]
  PIN m_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 57.840 680.000 58.440 ;
    END
  END m_in[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 676.000 6.840 680.000 7.440 ;
    END
  END rst
  PIN stall_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END stall_in
  PIN stall_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 4.000 ;
    END
  END stall_out
  PIN wishbone_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 676.000 2.210 680.000 ;
    END
  END wishbone_in[0]
  PIN wishbone_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 676.000 41.310 680.000 ;
    END
  END wishbone_in[10]
  PIN wishbone_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 676.000 44.990 680.000 ;
    END
  END wishbone_in[11]
  PIN wishbone_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 676.000 49.130 680.000 ;
    END
  END wishbone_in[12]
  PIN wishbone_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 676.000 53.270 680.000 ;
    END
  END wishbone_in[13]
  PIN wishbone_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 676.000 56.950 680.000 ;
    END
  END wishbone_in[14]
  PIN wishbone_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 676.000 61.090 680.000 ;
    END
  END wishbone_in[15]
  PIN wishbone_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 676.000 64.770 680.000 ;
    END
  END wishbone_in[16]
  PIN wishbone_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 676.000 68.910 680.000 ;
    END
  END wishbone_in[17]
  PIN wishbone_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 676.000 72.590 680.000 ;
    END
  END wishbone_in[18]
  PIN wishbone_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 676.000 76.730 680.000 ;
    END
  END wishbone_in[19]
  PIN wishbone_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 676.000 5.890 680.000 ;
    END
  END wishbone_in[1]
  PIN wishbone_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 676.000 80.410 680.000 ;
    END
  END wishbone_in[20]
  PIN wishbone_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 676.000 84.550 680.000 ;
    END
  END wishbone_in[21]
  PIN wishbone_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 676.000 88.230 680.000 ;
    END
  END wishbone_in[22]
  PIN wishbone_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 676.000 92.370 680.000 ;
    END
  END wishbone_in[23]
  PIN wishbone_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 676.000 96.510 680.000 ;
    END
  END wishbone_in[24]
  PIN wishbone_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 676.000 100.190 680.000 ;
    END
  END wishbone_in[25]
  PIN wishbone_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 676.000 104.330 680.000 ;
    END
  END wishbone_in[26]
  PIN wishbone_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 676.000 108.010 680.000 ;
    END
  END wishbone_in[27]
  PIN wishbone_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 676.000 112.150 680.000 ;
    END
  END wishbone_in[28]
  PIN wishbone_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 676.000 115.830 680.000 ;
    END
  END wishbone_in[29]
  PIN wishbone_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 676.000 10.030 680.000 ;
    END
  END wishbone_in[2]
  PIN wishbone_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 676.000 119.970 680.000 ;
    END
  END wishbone_in[30]
  PIN wishbone_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 676.000 123.650 680.000 ;
    END
  END wishbone_in[31]
  PIN wishbone_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 676.000 127.790 680.000 ;
    END
  END wishbone_in[32]
  PIN wishbone_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 676.000 131.470 680.000 ;
    END
  END wishbone_in[33]
  PIN wishbone_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 676.000 135.610 680.000 ;
    END
  END wishbone_in[34]
  PIN wishbone_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 676.000 139.750 680.000 ;
    END
  END wishbone_in[35]
  PIN wishbone_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 676.000 143.430 680.000 ;
    END
  END wishbone_in[36]
  PIN wishbone_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 676.000 147.570 680.000 ;
    END
  END wishbone_in[37]
  PIN wishbone_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 676.000 151.250 680.000 ;
    END
  END wishbone_in[38]
  PIN wishbone_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 676.000 155.390 680.000 ;
    END
  END wishbone_in[39]
  PIN wishbone_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 676.000 13.710 680.000 ;
    END
  END wishbone_in[3]
  PIN wishbone_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 676.000 159.070 680.000 ;
    END
  END wishbone_in[40]
  PIN wishbone_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 676.000 163.210 680.000 ;
    END
  END wishbone_in[41]
  PIN wishbone_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 676.000 166.890 680.000 ;
    END
  END wishbone_in[42]
  PIN wishbone_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 676.000 171.030 680.000 ;
    END
  END wishbone_in[43]
  PIN wishbone_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 676.000 174.710 680.000 ;
    END
  END wishbone_in[44]
  PIN wishbone_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 676.000 178.850 680.000 ;
    END
  END wishbone_in[45]
  PIN wishbone_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 676.000 182.530 680.000 ;
    END
  END wishbone_in[46]
  PIN wishbone_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 676.000 186.670 680.000 ;
    END
  END wishbone_in[47]
  PIN wishbone_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 676.000 190.810 680.000 ;
    END
  END wishbone_in[48]
  PIN wishbone_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 676.000 194.490 680.000 ;
    END
  END wishbone_in[49]
  PIN wishbone_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 676.000 17.850 680.000 ;
    END
  END wishbone_in[4]
  PIN wishbone_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 676.000 198.630 680.000 ;
    END
  END wishbone_in[50]
  PIN wishbone_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 676.000 202.310 680.000 ;
    END
  END wishbone_in[51]
  PIN wishbone_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 676.000 206.450 680.000 ;
    END
  END wishbone_in[52]
  PIN wishbone_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 676.000 210.130 680.000 ;
    END
  END wishbone_in[53]
  PIN wishbone_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 676.000 214.270 680.000 ;
    END
  END wishbone_in[54]
  PIN wishbone_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 676.000 217.950 680.000 ;
    END
  END wishbone_in[55]
  PIN wishbone_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 676.000 222.090 680.000 ;
    END
  END wishbone_in[56]
  PIN wishbone_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 676.000 225.770 680.000 ;
    END
  END wishbone_in[57]
  PIN wishbone_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 676.000 229.910 680.000 ;
    END
  END wishbone_in[58]
  PIN wishbone_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 676.000 234.050 680.000 ;
    END
  END wishbone_in[59]
  PIN wishbone_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 676.000 21.530 680.000 ;
    END
  END wishbone_in[5]
  PIN wishbone_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 676.000 237.730 680.000 ;
    END
  END wishbone_in[60]
  PIN wishbone_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 676.000 241.870 680.000 ;
    END
  END wishbone_in[61]
  PIN wishbone_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 676.000 245.550 680.000 ;
    END
  END wishbone_in[62]
  PIN wishbone_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 676.000 249.690 680.000 ;
    END
  END wishbone_in[63]
  PIN wishbone_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 676.000 253.370 680.000 ;
    END
  END wishbone_in[64]
  PIN wishbone_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 676.000 257.510 680.000 ;
    END
  END wishbone_in[65]
  PIN wishbone_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 676.000 25.670 680.000 ;
    END
  END wishbone_in[6]
  PIN wishbone_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 676.000 29.350 680.000 ;
    END
  END wishbone_in[7]
  PIN wishbone_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 676.000 33.490 680.000 ;
    END
  END wishbone_in[8]
  PIN wishbone_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 676.000 37.170 680.000 ;
    END
  END wishbone_in[9]
  PIN wishbone_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 676.000 261.190 680.000 ;
    END
  END wishbone_out[0]
  PIN wishbone_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 676.000 654.490 680.000 ;
    END
  END wishbone_out[100]
  PIN wishbone_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 676.000 658.170 680.000 ;
    END
  END wishbone_out[101]
  PIN wishbone_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 676.000 662.310 680.000 ;
    END
  END wishbone_out[102]
  PIN wishbone_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 676.000 665.990 680.000 ;
    END
  END wishbone_out[103]
  PIN wishbone_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 676.000 670.130 680.000 ;
    END
  END wishbone_out[104]
  PIN wishbone_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 676.000 673.810 680.000 ;
    END
  END wishbone_out[105]
  PIN wishbone_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 676.000 677.950 680.000 ;
    END
  END wishbone_out[106]
  PIN wishbone_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 676.000 300.750 680.000 ;
    END
  END wishbone_out[10]
  PIN wishbone_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 676.000 304.430 680.000 ;
    END
  END wishbone_out[11]
  PIN wishbone_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 676.000 308.570 680.000 ;
    END
  END wishbone_out[12]
  PIN wishbone_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 676.000 312.250 680.000 ;
    END
  END wishbone_out[13]
  PIN wishbone_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 676.000 316.390 680.000 ;
    END
  END wishbone_out[14]
  PIN wishbone_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 676.000 320.530 680.000 ;
    END
  END wishbone_out[15]
  PIN wishbone_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 676.000 324.210 680.000 ;
    END
  END wishbone_out[16]
  PIN wishbone_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 676.000 328.350 680.000 ;
    END
  END wishbone_out[17]
  PIN wishbone_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 676.000 332.030 680.000 ;
    END
  END wishbone_out[18]
  PIN wishbone_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 676.000 336.170 680.000 ;
    END
  END wishbone_out[19]
  PIN wishbone_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 676.000 265.330 680.000 ;
    END
  END wishbone_out[1]
  PIN wishbone_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 676.000 339.850 680.000 ;
    END
  END wishbone_out[20]
  PIN wishbone_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 676.000 343.990 680.000 ;
    END
  END wishbone_out[21]
  PIN wishbone_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 676.000 347.670 680.000 ;
    END
  END wishbone_out[22]
  PIN wishbone_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 676.000 351.810 680.000 ;
    END
  END wishbone_out[23]
  PIN wishbone_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 676.000 355.490 680.000 ;
    END
  END wishbone_out[24]
  PIN wishbone_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 676.000 359.630 680.000 ;
    END
  END wishbone_out[25]
  PIN wishbone_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 676.000 363.310 680.000 ;
    END
  END wishbone_out[26]
  PIN wishbone_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 676.000 367.450 680.000 ;
    END
  END wishbone_out[27]
  PIN wishbone_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 676.000 371.590 680.000 ;
    END
  END wishbone_out[28]
  PIN wishbone_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 676.000 375.270 680.000 ;
    END
  END wishbone_out[29]
  PIN wishbone_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 676.000 269.010 680.000 ;
    END
  END wishbone_out[2]
  PIN wishbone_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 676.000 379.410 680.000 ;
    END
  END wishbone_out[30]
  PIN wishbone_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 676.000 383.090 680.000 ;
    END
  END wishbone_out[31]
  PIN wishbone_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 676.000 387.230 680.000 ;
    END
  END wishbone_out[32]
  PIN wishbone_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 676.000 390.910 680.000 ;
    END
  END wishbone_out[33]
  PIN wishbone_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 676.000 395.050 680.000 ;
    END
  END wishbone_out[34]
  PIN wishbone_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 676.000 398.730 680.000 ;
    END
  END wishbone_out[35]
  PIN wishbone_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 676.000 402.870 680.000 ;
    END
  END wishbone_out[36]
  PIN wishbone_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 676.000 406.550 680.000 ;
    END
  END wishbone_out[37]
  PIN wishbone_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 676.000 410.690 680.000 ;
    END
  END wishbone_out[38]
  PIN wishbone_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 676.000 414.830 680.000 ;
    END
  END wishbone_out[39]
  PIN wishbone_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 676.000 273.150 680.000 ;
    END
  END wishbone_out[3]
  PIN wishbone_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 676.000 418.510 680.000 ;
    END
  END wishbone_out[40]
  PIN wishbone_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 676.000 422.650 680.000 ;
    END
  END wishbone_out[41]
  PIN wishbone_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 676.000 426.330 680.000 ;
    END
  END wishbone_out[42]
  PIN wishbone_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 676.000 430.470 680.000 ;
    END
  END wishbone_out[43]
  PIN wishbone_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 676.000 434.150 680.000 ;
    END
  END wishbone_out[44]
  PIN wishbone_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 676.000 438.290 680.000 ;
    END
  END wishbone_out[45]
  PIN wishbone_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 676.000 441.970 680.000 ;
    END
  END wishbone_out[46]
  PIN wishbone_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 676.000 446.110 680.000 ;
    END
  END wishbone_out[47]
  PIN wishbone_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 676.000 449.790 680.000 ;
    END
  END wishbone_out[48]
  PIN wishbone_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 676.000 453.930 680.000 ;
    END
  END wishbone_out[49]
  PIN wishbone_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 676.000 277.290 680.000 ;
    END
  END wishbone_out[4]
  PIN wishbone_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 676.000 458.070 680.000 ;
    END
  END wishbone_out[50]
  PIN wishbone_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 676.000 461.750 680.000 ;
    END
  END wishbone_out[51]
  PIN wishbone_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 676.000 465.890 680.000 ;
    END
  END wishbone_out[52]
  PIN wishbone_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 676.000 469.570 680.000 ;
    END
  END wishbone_out[53]
  PIN wishbone_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 676.000 473.710 680.000 ;
    END
  END wishbone_out[54]
  PIN wishbone_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 676.000 477.390 680.000 ;
    END
  END wishbone_out[55]
  PIN wishbone_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 676.000 481.530 680.000 ;
    END
  END wishbone_out[56]
  PIN wishbone_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 676.000 485.210 680.000 ;
    END
  END wishbone_out[57]
  PIN wishbone_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 676.000 489.350 680.000 ;
    END
  END wishbone_out[58]
  PIN wishbone_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 676.000 493.030 680.000 ;
    END
  END wishbone_out[59]
  PIN wishbone_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 676.000 280.970 680.000 ;
    END
  END wishbone_out[5]
  PIN wishbone_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 676.000 497.170 680.000 ;
    END
  END wishbone_out[60]
  PIN wishbone_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 676.000 501.310 680.000 ;
    END
  END wishbone_out[61]
  PIN wishbone_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 676.000 504.990 680.000 ;
    END
  END wishbone_out[62]
  PIN wishbone_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 676.000 509.130 680.000 ;
    END
  END wishbone_out[63]
  PIN wishbone_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 676.000 512.810 680.000 ;
    END
  END wishbone_out[64]
  PIN wishbone_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 676.000 516.950 680.000 ;
    END
  END wishbone_out[65]
  PIN wishbone_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 676.000 520.630 680.000 ;
    END
  END wishbone_out[66]
  PIN wishbone_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 676.000 524.770 680.000 ;
    END
  END wishbone_out[67]
  PIN wishbone_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 676.000 528.450 680.000 ;
    END
  END wishbone_out[68]
  PIN wishbone_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 676.000 532.590 680.000 ;
    END
  END wishbone_out[69]
  PIN wishbone_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 676.000 285.110 680.000 ;
    END
  END wishbone_out[6]
  PIN wishbone_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 676.000 536.270 680.000 ;
    END
  END wishbone_out[70]
  PIN wishbone_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 676.000 540.410 680.000 ;
    END
  END wishbone_out[71]
  PIN wishbone_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 676.000 544.090 680.000 ;
    END
  END wishbone_out[72]
  PIN wishbone_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 676.000 548.230 680.000 ;
    END
  END wishbone_out[73]
  PIN wishbone_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 676.000 552.370 680.000 ;
    END
  END wishbone_out[74]
  PIN wishbone_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 676.000 556.050 680.000 ;
    END
  END wishbone_out[75]
  PIN wishbone_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 676.000 560.190 680.000 ;
    END
  END wishbone_out[76]
  PIN wishbone_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 676.000 563.870 680.000 ;
    END
  END wishbone_out[77]
  PIN wishbone_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 676.000 568.010 680.000 ;
    END
  END wishbone_out[78]
  PIN wishbone_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 676.000 571.690 680.000 ;
    END
  END wishbone_out[79]
  PIN wishbone_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 676.000 288.790 680.000 ;
    END
  END wishbone_out[7]
  PIN wishbone_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 676.000 575.830 680.000 ;
    END
  END wishbone_out[80]
  PIN wishbone_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 676.000 579.510 680.000 ;
    END
  END wishbone_out[81]
  PIN wishbone_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 676.000 583.650 680.000 ;
    END
  END wishbone_out[82]
  PIN wishbone_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 676.000 587.330 680.000 ;
    END
  END wishbone_out[83]
  PIN wishbone_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 676.000 591.470 680.000 ;
    END
  END wishbone_out[84]
  PIN wishbone_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 676.000 595.610 680.000 ;
    END
  END wishbone_out[85]
  PIN wishbone_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 676.000 599.290 680.000 ;
    END
  END wishbone_out[86]
  PIN wishbone_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 676.000 603.430 680.000 ;
    END
  END wishbone_out[87]
  PIN wishbone_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 676.000 607.110 680.000 ;
    END
  END wishbone_out[88]
  PIN wishbone_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 676.000 611.250 680.000 ;
    END
  END wishbone_out[89]
  PIN wishbone_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 676.000 292.930 680.000 ;
    END
  END wishbone_out[8]
  PIN wishbone_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 676.000 614.930 680.000 ;
    END
  END wishbone_out[90]
  PIN wishbone_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 676.000 619.070 680.000 ;
    END
  END wishbone_out[91]
  PIN wishbone_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 676.000 622.750 680.000 ;
    END
  END wishbone_out[92]
  PIN wishbone_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 676.000 626.890 680.000 ;
    END
  END wishbone_out[93]
  PIN wishbone_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 676.000 630.570 680.000 ;
    END
  END wishbone_out[94]
  PIN wishbone_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 676.000 634.710 680.000 ;
    END
  END wishbone_out[95]
  PIN wishbone_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 676.000 638.850 680.000 ;
    END
  END wishbone_out[96]
  PIN wishbone_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 676.000 642.530 680.000 ;
    END
  END wishbone_out[97]
  PIN wishbone_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 676.000 646.670 680.000 ;
    END
  END wishbone_out[98]
  PIN wishbone_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 676.000 650.350 680.000 ;
    END
  END wishbone_out[99]
  PIN wishbone_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 676.000 296.610 680.000 ;
    END
  END wishbone_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 669.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 669.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 669.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 669.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 669.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 669.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 669.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 669.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 669.360 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 674.360 669.205 ;
      LAYER met1 ;
        RECT 1.910 0.040 677.970 669.760 ;
      LAYER met2 ;
        RECT 2.490 675.720 5.330 676.000 ;
        RECT 6.170 675.720 9.470 676.000 ;
        RECT 10.310 675.720 13.150 676.000 ;
        RECT 13.990 675.720 17.290 676.000 ;
        RECT 18.130 675.720 20.970 676.000 ;
        RECT 21.810 675.720 25.110 676.000 ;
        RECT 25.950 675.720 28.790 676.000 ;
        RECT 29.630 675.720 32.930 676.000 ;
        RECT 33.770 675.720 36.610 676.000 ;
        RECT 37.450 675.720 40.750 676.000 ;
        RECT 41.590 675.720 44.430 676.000 ;
        RECT 45.270 675.720 48.570 676.000 ;
        RECT 49.410 675.720 52.710 676.000 ;
        RECT 53.550 675.720 56.390 676.000 ;
        RECT 57.230 675.720 60.530 676.000 ;
        RECT 61.370 675.720 64.210 676.000 ;
        RECT 65.050 675.720 68.350 676.000 ;
        RECT 69.190 675.720 72.030 676.000 ;
        RECT 72.870 675.720 76.170 676.000 ;
        RECT 77.010 675.720 79.850 676.000 ;
        RECT 80.690 675.720 83.990 676.000 ;
        RECT 84.830 675.720 87.670 676.000 ;
        RECT 88.510 675.720 91.810 676.000 ;
        RECT 92.650 675.720 95.950 676.000 ;
        RECT 96.790 675.720 99.630 676.000 ;
        RECT 100.470 675.720 103.770 676.000 ;
        RECT 104.610 675.720 107.450 676.000 ;
        RECT 108.290 675.720 111.590 676.000 ;
        RECT 112.430 675.720 115.270 676.000 ;
        RECT 116.110 675.720 119.410 676.000 ;
        RECT 120.250 675.720 123.090 676.000 ;
        RECT 123.930 675.720 127.230 676.000 ;
        RECT 128.070 675.720 130.910 676.000 ;
        RECT 131.750 675.720 135.050 676.000 ;
        RECT 135.890 675.720 139.190 676.000 ;
        RECT 140.030 675.720 142.870 676.000 ;
        RECT 143.710 675.720 147.010 676.000 ;
        RECT 147.850 675.720 150.690 676.000 ;
        RECT 151.530 675.720 154.830 676.000 ;
        RECT 155.670 675.720 158.510 676.000 ;
        RECT 159.350 675.720 162.650 676.000 ;
        RECT 163.490 675.720 166.330 676.000 ;
        RECT 167.170 675.720 170.470 676.000 ;
        RECT 171.310 675.720 174.150 676.000 ;
        RECT 174.990 675.720 178.290 676.000 ;
        RECT 179.130 675.720 181.970 676.000 ;
        RECT 182.810 675.720 186.110 676.000 ;
        RECT 186.950 675.720 190.250 676.000 ;
        RECT 191.090 675.720 193.930 676.000 ;
        RECT 194.770 675.720 198.070 676.000 ;
        RECT 198.910 675.720 201.750 676.000 ;
        RECT 202.590 675.720 205.890 676.000 ;
        RECT 206.730 675.720 209.570 676.000 ;
        RECT 210.410 675.720 213.710 676.000 ;
        RECT 214.550 675.720 217.390 676.000 ;
        RECT 218.230 675.720 221.530 676.000 ;
        RECT 222.370 675.720 225.210 676.000 ;
        RECT 226.050 675.720 229.350 676.000 ;
        RECT 230.190 675.720 233.490 676.000 ;
        RECT 234.330 675.720 237.170 676.000 ;
        RECT 238.010 675.720 241.310 676.000 ;
        RECT 242.150 675.720 244.990 676.000 ;
        RECT 245.830 675.720 249.130 676.000 ;
        RECT 249.970 675.720 252.810 676.000 ;
        RECT 253.650 675.720 256.950 676.000 ;
        RECT 257.790 675.720 260.630 676.000 ;
        RECT 261.470 675.720 264.770 676.000 ;
        RECT 265.610 675.720 268.450 676.000 ;
        RECT 269.290 675.720 272.590 676.000 ;
        RECT 273.430 675.720 276.730 676.000 ;
        RECT 277.570 675.720 280.410 676.000 ;
        RECT 281.250 675.720 284.550 676.000 ;
        RECT 285.390 675.720 288.230 676.000 ;
        RECT 289.070 675.720 292.370 676.000 ;
        RECT 293.210 675.720 296.050 676.000 ;
        RECT 296.890 675.720 300.190 676.000 ;
        RECT 301.030 675.720 303.870 676.000 ;
        RECT 304.710 675.720 308.010 676.000 ;
        RECT 308.850 675.720 311.690 676.000 ;
        RECT 312.530 675.720 315.830 676.000 ;
        RECT 316.670 675.720 319.970 676.000 ;
        RECT 320.810 675.720 323.650 676.000 ;
        RECT 324.490 675.720 327.790 676.000 ;
        RECT 328.630 675.720 331.470 676.000 ;
        RECT 332.310 675.720 335.610 676.000 ;
        RECT 336.450 675.720 339.290 676.000 ;
        RECT 340.130 675.720 343.430 676.000 ;
        RECT 344.270 675.720 347.110 676.000 ;
        RECT 347.950 675.720 351.250 676.000 ;
        RECT 352.090 675.720 354.930 676.000 ;
        RECT 355.770 675.720 359.070 676.000 ;
        RECT 359.910 675.720 362.750 676.000 ;
        RECT 363.590 675.720 366.890 676.000 ;
        RECT 367.730 675.720 371.030 676.000 ;
        RECT 371.870 675.720 374.710 676.000 ;
        RECT 375.550 675.720 378.850 676.000 ;
        RECT 379.690 675.720 382.530 676.000 ;
        RECT 383.370 675.720 386.670 676.000 ;
        RECT 387.510 675.720 390.350 676.000 ;
        RECT 391.190 675.720 394.490 676.000 ;
        RECT 395.330 675.720 398.170 676.000 ;
        RECT 399.010 675.720 402.310 676.000 ;
        RECT 403.150 675.720 405.990 676.000 ;
        RECT 406.830 675.720 410.130 676.000 ;
        RECT 410.970 675.720 414.270 676.000 ;
        RECT 415.110 675.720 417.950 676.000 ;
        RECT 418.790 675.720 422.090 676.000 ;
        RECT 422.930 675.720 425.770 676.000 ;
        RECT 426.610 675.720 429.910 676.000 ;
        RECT 430.750 675.720 433.590 676.000 ;
        RECT 434.430 675.720 437.730 676.000 ;
        RECT 438.570 675.720 441.410 676.000 ;
        RECT 442.250 675.720 445.550 676.000 ;
        RECT 446.390 675.720 449.230 676.000 ;
        RECT 450.070 675.720 453.370 676.000 ;
        RECT 454.210 675.720 457.510 676.000 ;
        RECT 458.350 675.720 461.190 676.000 ;
        RECT 462.030 675.720 465.330 676.000 ;
        RECT 466.170 675.720 469.010 676.000 ;
        RECT 469.850 675.720 473.150 676.000 ;
        RECT 473.990 675.720 476.830 676.000 ;
        RECT 477.670 675.720 480.970 676.000 ;
        RECT 481.810 675.720 484.650 676.000 ;
        RECT 485.490 675.720 488.790 676.000 ;
        RECT 489.630 675.720 492.470 676.000 ;
        RECT 493.310 675.720 496.610 676.000 ;
        RECT 497.450 675.720 500.750 676.000 ;
        RECT 501.590 675.720 504.430 676.000 ;
        RECT 505.270 675.720 508.570 676.000 ;
        RECT 509.410 675.720 512.250 676.000 ;
        RECT 513.090 675.720 516.390 676.000 ;
        RECT 517.230 675.720 520.070 676.000 ;
        RECT 520.910 675.720 524.210 676.000 ;
        RECT 525.050 675.720 527.890 676.000 ;
        RECT 528.730 675.720 532.030 676.000 ;
        RECT 532.870 675.720 535.710 676.000 ;
        RECT 536.550 675.720 539.850 676.000 ;
        RECT 540.690 675.720 543.530 676.000 ;
        RECT 544.370 675.720 547.670 676.000 ;
        RECT 548.510 675.720 551.810 676.000 ;
        RECT 552.650 675.720 555.490 676.000 ;
        RECT 556.330 675.720 559.630 676.000 ;
        RECT 560.470 675.720 563.310 676.000 ;
        RECT 564.150 675.720 567.450 676.000 ;
        RECT 568.290 675.720 571.130 676.000 ;
        RECT 571.970 675.720 575.270 676.000 ;
        RECT 576.110 675.720 578.950 676.000 ;
        RECT 579.790 675.720 583.090 676.000 ;
        RECT 583.930 675.720 586.770 676.000 ;
        RECT 587.610 675.720 590.910 676.000 ;
        RECT 591.750 675.720 595.050 676.000 ;
        RECT 595.890 675.720 598.730 676.000 ;
        RECT 599.570 675.720 602.870 676.000 ;
        RECT 603.710 675.720 606.550 676.000 ;
        RECT 607.390 675.720 610.690 676.000 ;
        RECT 611.530 675.720 614.370 676.000 ;
        RECT 615.210 675.720 618.510 676.000 ;
        RECT 619.350 675.720 622.190 676.000 ;
        RECT 623.030 675.720 626.330 676.000 ;
        RECT 627.170 675.720 630.010 676.000 ;
        RECT 630.850 675.720 634.150 676.000 ;
        RECT 634.990 675.720 638.290 676.000 ;
        RECT 639.130 675.720 641.970 676.000 ;
        RECT 642.810 675.720 646.110 676.000 ;
        RECT 646.950 675.720 649.790 676.000 ;
        RECT 650.630 675.720 653.930 676.000 ;
        RECT 654.770 675.720 657.610 676.000 ;
        RECT 658.450 675.720 661.750 676.000 ;
        RECT 662.590 675.720 665.430 676.000 ;
        RECT 666.270 675.720 669.570 676.000 ;
        RECT 670.410 675.720 673.250 676.000 ;
        RECT 674.090 675.720 677.390 676.000 ;
        RECT 1.940 4.280 677.940 675.720 ;
        RECT 2.490 0.010 5.330 4.280 ;
        RECT 6.170 0.010 9.470 4.280 ;
        RECT 10.310 0.010 13.150 4.280 ;
        RECT 13.990 0.010 17.290 4.280 ;
        RECT 18.130 0.010 20.970 4.280 ;
        RECT 21.810 0.010 25.110 4.280 ;
        RECT 25.950 0.010 28.790 4.280 ;
        RECT 29.630 0.010 32.930 4.280 ;
        RECT 33.770 0.010 36.610 4.280 ;
        RECT 37.450 0.010 40.750 4.280 ;
        RECT 41.590 0.010 44.430 4.280 ;
        RECT 45.270 0.010 48.570 4.280 ;
        RECT 49.410 0.010 52.710 4.280 ;
        RECT 53.550 0.010 56.390 4.280 ;
        RECT 57.230 0.010 60.530 4.280 ;
        RECT 61.370 0.010 64.210 4.280 ;
        RECT 65.050 0.010 68.350 4.280 ;
        RECT 69.190 0.010 72.030 4.280 ;
        RECT 72.870 0.010 76.170 4.280 ;
        RECT 77.010 0.010 79.850 4.280 ;
        RECT 80.690 0.010 83.990 4.280 ;
        RECT 84.830 0.010 87.670 4.280 ;
        RECT 88.510 0.010 91.810 4.280 ;
        RECT 92.650 0.010 95.950 4.280 ;
        RECT 96.790 0.010 99.630 4.280 ;
        RECT 100.470 0.010 103.770 4.280 ;
        RECT 104.610 0.010 107.450 4.280 ;
        RECT 108.290 0.010 111.590 4.280 ;
        RECT 112.430 0.010 115.270 4.280 ;
        RECT 116.110 0.010 119.410 4.280 ;
        RECT 120.250 0.010 123.090 4.280 ;
        RECT 123.930 0.010 127.230 4.280 ;
        RECT 128.070 0.010 130.910 4.280 ;
        RECT 131.750 0.010 135.050 4.280 ;
        RECT 135.890 0.010 139.190 4.280 ;
        RECT 140.030 0.010 142.870 4.280 ;
        RECT 143.710 0.010 147.010 4.280 ;
        RECT 147.850 0.010 150.690 4.280 ;
        RECT 151.530 0.010 154.830 4.280 ;
        RECT 155.670 0.010 158.510 4.280 ;
        RECT 159.350 0.010 162.650 4.280 ;
        RECT 163.490 0.010 166.330 4.280 ;
        RECT 167.170 0.010 170.470 4.280 ;
        RECT 171.310 0.010 174.150 4.280 ;
        RECT 174.990 0.010 178.290 4.280 ;
        RECT 179.130 0.010 181.970 4.280 ;
        RECT 182.810 0.010 186.110 4.280 ;
        RECT 186.950 0.010 190.250 4.280 ;
        RECT 191.090 0.010 193.930 4.280 ;
        RECT 194.770 0.010 198.070 4.280 ;
        RECT 198.910 0.010 201.750 4.280 ;
        RECT 202.590 0.010 205.890 4.280 ;
        RECT 206.730 0.010 209.570 4.280 ;
        RECT 210.410 0.010 213.710 4.280 ;
        RECT 214.550 0.010 217.390 4.280 ;
        RECT 218.230 0.010 221.530 4.280 ;
        RECT 222.370 0.010 225.210 4.280 ;
        RECT 226.050 0.010 229.350 4.280 ;
        RECT 230.190 0.010 233.490 4.280 ;
        RECT 234.330 0.010 237.170 4.280 ;
        RECT 238.010 0.010 241.310 4.280 ;
        RECT 242.150 0.010 244.990 4.280 ;
        RECT 245.830 0.010 249.130 4.280 ;
        RECT 249.970 0.010 252.810 4.280 ;
        RECT 253.650 0.010 256.950 4.280 ;
        RECT 257.790 0.010 260.630 4.280 ;
        RECT 261.470 0.010 264.770 4.280 ;
        RECT 265.610 0.010 268.450 4.280 ;
        RECT 269.290 0.010 272.590 4.280 ;
        RECT 273.430 0.010 276.730 4.280 ;
        RECT 277.570 0.010 280.410 4.280 ;
        RECT 281.250 0.010 284.550 4.280 ;
        RECT 285.390 0.010 288.230 4.280 ;
        RECT 289.070 0.010 292.370 4.280 ;
        RECT 293.210 0.010 296.050 4.280 ;
        RECT 296.890 0.010 300.190 4.280 ;
        RECT 301.030 0.010 303.870 4.280 ;
        RECT 304.710 0.010 308.010 4.280 ;
        RECT 308.850 0.010 311.690 4.280 ;
        RECT 312.530 0.010 315.830 4.280 ;
        RECT 316.670 0.010 319.970 4.280 ;
        RECT 320.810 0.010 323.650 4.280 ;
        RECT 324.490 0.010 327.790 4.280 ;
        RECT 328.630 0.010 331.470 4.280 ;
        RECT 332.310 0.010 335.610 4.280 ;
        RECT 336.450 0.010 339.290 4.280 ;
        RECT 340.130 0.010 343.430 4.280 ;
        RECT 344.270 0.010 347.110 4.280 ;
        RECT 347.950 0.010 351.250 4.280 ;
        RECT 352.090 0.010 354.930 4.280 ;
        RECT 355.770 0.010 359.070 4.280 ;
        RECT 359.910 0.010 362.750 4.280 ;
        RECT 363.590 0.010 366.890 4.280 ;
        RECT 367.730 0.010 371.030 4.280 ;
        RECT 371.870 0.010 374.710 4.280 ;
        RECT 375.550 0.010 378.850 4.280 ;
        RECT 379.690 0.010 382.530 4.280 ;
        RECT 383.370 0.010 386.670 4.280 ;
        RECT 387.510 0.010 390.350 4.280 ;
        RECT 391.190 0.010 394.490 4.280 ;
        RECT 395.330 0.010 398.170 4.280 ;
        RECT 399.010 0.010 402.310 4.280 ;
        RECT 403.150 0.010 405.990 4.280 ;
        RECT 406.830 0.010 410.130 4.280 ;
        RECT 410.970 0.010 414.270 4.280 ;
        RECT 415.110 0.010 417.950 4.280 ;
        RECT 418.790 0.010 422.090 4.280 ;
        RECT 422.930 0.010 425.770 4.280 ;
        RECT 426.610 0.010 429.910 4.280 ;
        RECT 430.750 0.010 433.590 4.280 ;
        RECT 434.430 0.010 437.730 4.280 ;
        RECT 438.570 0.010 441.410 4.280 ;
        RECT 442.250 0.010 445.550 4.280 ;
        RECT 446.390 0.010 449.230 4.280 ;
        RECT 450.070 0.010 453.370 4.280 ;
        RECT 454.210 0.010 457.510 4.280 ;
        RECT 458.350 0.010 461.190 4.280 ;
        RECT 462.030 0.010 465.330 4.280 ;
        RECT 466.170 0.010 469.010 4.280 ;
        RECT 469.850 0.010 473.150 4.280 ;
        RECT 473.990 0.010 476.830 4.280 ;
        RECT 477.670 0.010 480.970 4.280 ;
        RECT 481.810 0.010 484.650 4.280 ;
        RECT 485.490 0.010 488.790 4.280 ;
        RECT 489.630 0.010 492.470 4.280 ;
        RECT 493.310 0.010 496.610 4.280 ;
        RECT 497.450 0.010 500.750 4.280 ;
        RECT 501.590 0.010 504.430 4.280 ;
        RECT 505.270 0.010 508.570 4.280 ;
        RECT 509.410 0.010 512.250 4.280 ;
        RECT 513.090 0.010 516.390 4.280 ;
        RECT 517.230 0.010 520.070 4.280 ;
        RECT 520.910 0.010 524.210 4.280 ;
        RECT 525.050 0.010 527.890 4.280 ;
        RECT 528.730 0.010 532.030 4.280 ;
        RECT 532.870 0.010 535.710 4.280 ;
        RECT 536.550 0.010 539.850 4.280 ;
        RECT 540.690 0.010 543.530 4.280 ;
        RECT 544.370 0.010 547.670 4.280 ;
        RECT 548.510 0.010 551.810 4.280 ;
        RECT 552.650 0.010 555.490 4.280 ;
        RECT 556.330 0.010 559.630 4.280 ;
        RECT 560.470 0.010 563.310 4.280 ;
        RECT 564.150 0.010 567.450 4.280 ;
        RECT 568.290 0.010 571.130 4.280 ;
        RECT 571.970 0.010 575.270 4.280 ;
        RECT 576.110 0.010 578.950 4.280 ;
        RECT 579.790 0.010 583.090 4.280 ;
        RECT 583.930 0.010 586.770 4.280 ;
        RECT 587.610 0.010 590.910 4.280 ;
        RECT 591.750 0.010 595.050 4.280 ;
        RECT 595.890 0.010 598.730 4.280 ;
        RECT 599.570 0.010 602.870 4.280 ;
        RECT 603.710 0.010 606.550 4.280 ;
        RECT 607.390 0.010 610.690 4.280 ;
        RECT 611.530 0.010 614.370 4.280 ;
        RECT 615.210 0.010 618.510 4.280 ;
        RECT 619.350 0.010 622.190 4.280 ;
        RECT 623.030 0.010 626.330 4.280 ;
        RECT 627.170 0.010 630.010 4.280 ;
        RECT 630.850 0.010 634.150 4.280 ;
        RECT 634.990 0.010 638.290 4.280 ;
        RECT 639.130 0.010 641.970 4.280 ;
        RECT 642.810 0.010 646.110 4.280 ;
        RECT 646.950 0.010 649.790 4.280 ;
        RECT 650.630 0.010 653.930 4.280 ;
        RECT 654.770 0.010 657.610 4.280 ;
        RECT 658.450 0.010 661.750 4.280 ;
        RECT 662.590 0.010 665.430 4.280 ;
        RECT 666.270 0.010 669.570 4.280 ;
        RECT 670.410 0.010 673.250 4.280 ;
        RECT 674.090 0.010 677.390 4.280 ;
      LAYER met3 ;
        RECT 14.325 667.440 676.000 669.285 ;
        RECT 14.325 666.040 675.600 667.440 ;
        RECT 14.325 662.000 676.000 666.040 ;
        RECT 14.325 660.600 675.600 662.000 ;
        RECT 14.325 657.240 676.000 660.600 ;
        RECT 14.325 655.840 675.600 657.240 ;
        RECT 14.325 651.800 676.000 655.840 ;
        RECT 14.325 650.400 675.600 651.800 ;
        RECT 14.325 647.040 676.000 650.400 ;
        RECT 14.325 645.640 675.600 647.040 ;
        RECT 14.325 641.600 676.000 645.640 ;
        RECT 14.325 640.200 675.600 641.600 ;
        RECT 14.325 636.840 676.000 640.200 ;
        RECT 14.325 635.440 675.600 636.840 ;
        RECT 14.325 631.400 676.000 635.440 ;
        RECT 14.325 630.000 675.600 631.400 ;
        RECT 14.325 626.640 676.000 630.000 ;
        RECT 14.325 625.240 675.600 626.640 ;
        RECT 14.325 621.200 676.000 625.240 ;
        RECT 14.325 619.800 675.600 621.200 ;
        RECT 14.325 616.440 676.000 619.800 ;
        RECT 14.325 615.040 675.600 616.440 ;
        RECT 14.325 611.000 676.000 615.040 ;
        RECT 14.325 609.600 675.600 611.000 ;
        RECT 14.325 606.240 676.000 609.600 ;
        RECT 14.325 604.840 675.600 606.240 ;
        RECT 14.325 600.800 676.000 604.840 ;
        RECT 14.325 599.400 675.600 600.800 ;
        RECT 14.325 596.040 676.000 599.400 ;
        RECT 14.325 594.640 675.600 596.040 ;
        RECT 14.325 590.600 676.000 594.640 ;
        RECT 14.325 589.200 675.600 590.600 ;
        RECT 14.325 585.840 676.000 589.200 ;
        RECT 14.325 584.440 675.600 585.840 ;
        RECT 14.325 580.400 676.000 584.440 ;
        RECT 14.325 579.000 675.600 580.400 ;
        RECT 14.325 575.640 676.000 579.000 ;
        RECT 14.325 574.240 675.600 575.640 ;
        RECT 14.325 570.200 676.000 574.240 ;
        RECT 14.325 568.800 675.600 570.200 ;
        RECT 14.325 565.440 676.000 568.800 ;
        RECT 14.325 564.040 675.600 565.440 ;
        RECT 14.325 560.000 676.000 564.040 ;
        RECT 14.325 558.600 675.600 560.000 ;
        RECT 14.325 555.240 676.000 558.600 ;
        RECT 14.325 553.840 675.600 555.240 ;
        RECT 14.325 549.800 676.000 553.840 ;
        RECT 14.325 548.400 675.600 549.800 ;
        RECT 14.325 544.360 676.000 548.400 ;
        RECT 14.325 542.960 675.600 544.360 ;
        RECT 14.325 539.600 676.000 542.960 ;
        RECT 14.325 538.200 675.600 539.600 ;
        RECT 14.325 534.160 676.000 538.200 ;
        RECT 14.325 532.760 675.600 534.160 ;
        RECT 14.325 529.400 676.000 532.760 ;
        RECT 14.325 528.000 675.600 529.400 ;
        RECT 14.325 523.960 676.000 528.000 ;
        RECT 14.325 522.560 675.600 523.960 ;
        RECT 14.325 519.200 676.000 522.560 ;
        RECT 14.325 517.800 675.600 519.200 ;
        RECT 14.325 513.760 676.000 517.800 ;
        RECT 14.325 512.360 675.600 513.760 ;
        RECT 14.325 509.000 676.000 512.360 ;
        RECT 14.325 507.600 675.600 509.000 ;
        RECT 14.325 503.560 676.000 507.600 ;
        RECT 14.325 502.160 675.600 503.560 ;
        RECT 14.325 498.800 676.000 502.160 ;
        RECT 14.325 497.400 675.600 498.800 ;
        RECT 14.325 493.360 676.000 497.400 ;
        RECT 14.325 491.960 675.600 493.360 ;
        RECT 14.325 488.600 676.000 491.960 ;
        RECT 14.325 487.200 675.600 488.600 ;
        RECT 14.325 483.160 676.000 487.200 ;
        RECT 14.325 481.760 675.600 483.160 ;
        RECT 14.325 478.400 676.000 481.760 ;
        RECT 14.325 477.000 675.600 478.400 ;
        RECT 14.325 472.960 676.000 477.000 ;
        RECT 14.325 471.560 675.600 472.960 ;
        RECT 14.325 468.200 676.000 471.560 ;
        RECT 14.325 466.800 675.600 468.200 ;
        RECT 14.325 462.760 676.000 466.800 ;
        RECT 14.325 461.360 675.600 462.760 ;
        RECT 14.325 458.000 676.000 461.360 ;
        RECT 14.325 456.600 675.600 458.000 ;
        RECT 14.325 452.560 676.000 456.600 ;
        RECT 14.325 451.160 675.600 452.560 ;
        RECT 14.325 447.800 676.000 451.160 ;
        RECT 14.325 446.400 675.600 447.800 ;
        RECT 14.325 442.360 676.000 446.400 ;
        RECT 14.325 440.960 675.600 442.360 ;
        RECT 14.325 437.600 676.000 440.960 ;
        RECT 14.325 436.200 675.600 437.600 ;
        RECT 14.325 432.160 676.000 436.200 ;
        RECT 14.325 430.760 675.600 432.160 ;
        RECT 14.325 427.400 676.000 430.760 ;
        RECT 14.325 426.000 675.600 427.400 ;
        RECT 14.325 421.960 676.000 426.000 ;
        RECT 14.325 420.560 675.600 421.960 ;
        RECT 14.325 417.200 676.000 420.560 ;
        RECT 14.325 415.800 675.600 417.200 ;
        RECT 14.325 411.760 676.000 415.800 ;
        RECT 14.325 410.360 675.600 411.760 ;
        RECT 14.325 406.320 676.000 410.360 ;
        RECT 14.325 404.920 675.600 406.320 ;
        RECT 14.325 401.560 676.000 404.920 ;
        RECT 14.325 400.160 675.600 401.560 ;
        RECT 14.325 396.120 676.000 400.160 ;
        RECT 14.325 394.720 675.600 396.120 ;
        RECT 14.325 391.360 676.000 394.720 ;
        RECT 14.325 389.960 675.600 391.360 ;
        RECT 14.325 385.920 676.000 389.960 ;
        RECT 14.325 384.520 675.600 385.920 ;
        RECT 14.325 381.160 676.000 384.520 ;
        RECT 14.325 379.760 675.600 381.160 ;
        RECT 14.325 375.720 676.000 379.760 ;
        RECT 14.325 374.320 675.600 375.720 ;
        RECT 14.325 370.960 676.000 374.320 ;
        RECT 14.325 369.560 675.600 370.960 ;
        RECT 14.325 365.520 676.000 369.560 ;
        RECT 14.325 364.120 675.600 365.520 ;
        RECT 14.325 360.760 676.000 364.120 ;
        RECT 14.325 359.360 675.600 360.760 ;
        RECT 14.325 355.320 676.000 359.360 ;
        RECT 14.325 353.920 675.600 355.320 ;
        RECT 14.325 350.560 676.000 353.920 ;
        RECT 14.325 349.160 675.600 350.560 ;
        RECT 14.325 345.120 676.000 349.160 ;
        RECT 14.325 343.720 675.600 345.120 ;
        RECT 14.325 340.360 676.000 343.720 ;
        RECT 14.325 338.960 675.600 340.360 ;
        RECT 14.325 334.920 676.000 338.960 ;
        RECT 14.325 333.520 675.600 334.920 ;
        RECT 14.325 330.160 676.000 333.520 ;
        RECT 14.325 328.760 675.600 330.160 ;
        RECT 14.325 324.720 676.000 328.760 ;
        RECT 14.325 323.320 675.600 324.720 ;
        RECT 14.325 319.960 676.000 323.320 ;
        RECT 14.325 318.560 675.600 319.960 ;
        RECT 14.325 314.520 676.000 318.560 ;
        RECT 14.325 313.120 675.600 314.520 ;
        RECT 14.325 309.760 676.000 313.120 ;
        RECT 14.325 308.360 675.600 309.760 ;
        RECT 14.325 304.320 676.000 308.360 ;
        RECT 14.325 302.920 675.600 304.320 ;
        RECT 14.325 299.560 676.000 302.920 ;
        RECT 14.325 298.160 675.600 299.560 ;
        RECT 14.325 294.120 676.000 298.160 ;
        RECT 14.325 292.720 675.600 294.120 ;
        RECT 14.325 289.360 676.000 292.720 ;
        RECT 14.325 287.960 675.600 289.360 ;
        RECT 14.325 283.920 676.000 287.960 ;
        RECT 14.325 282.520 675.600 283.920 ;
        RECT 14.325 279.160 676.000 282.520 ;
        RECT 14.325 277.760 675.600 279.160 ;
        RECT 14.325 273.720 676.000 277.760 ;
        RECT 14.325 272.320 675.600 273.720 ;
        RECT 14.325 268.280 676.000 272.320 ;
        RECT 14.325 266.880 675.600 268.280 ;
        RECT 14.325 263.520 676.000 266.880 ;
        RECT 14.325 262.120 675.600 263.520 ;
        RECT 14.325 258.080 676.000 262.120 ;
        RECT 14.325 256.680 675.600 258.080 ;
        RECT 14.325 253.320 676.000 256.680 ;
        RECT 14.325 251.920 675.600 253.320 ;
        RECT 14.325 247.880 676.000 251.920 ;
        RECT 14.325 246.480 675.600 247.880 ;
        RECT 14.325 243.120 676.000 246.480 ;
        RECT 14.325 241.720 675.600 243.120 ;
        RECT 14.325 237.680 676.000 241.720 ;
        RECT 14.325 236.280 675.600 237.680 ;
        RECT 14.325 232.920 676.000 236.280 ;
        RECT 14.325 231.520 675.600 232.920 ;
        RECT 14.325 227.480 676.000 231.520 ;
        RECT 14.325 226.080 675.600 227.480 ;
        RECT 14.325 222.720 676.000 226.080 ;
        RECT 14.325 221.320 675.600 222.720 ;
        RECT 14.325 217.280 676.000 221.320 ;
        RECT 14.325 215.880 675.600 217.280 ;
        RECT 14.325 212.520 676.000 215.880 ;
        RECT 14.325 211.120 675.600 212.520 ;
        RECT 14.325 207.080 676.000 211.120 ;
        RECT 14.325 205.680 675.600 207.080 ;
        RECT 14.325 202.320 676.000 205.680 ;
        RECT 14.325 200.920 675.600 202.320 ;
        RECT 14.325 196.880 676.000 200.920 ;
        RECT 14.325 195.480 675.600 196.880 ;
        RECT 14.325 192.120 676.000 195.480 ;
        RECT 14.325 190.720 675.600 192.120 ;
        RECT 14.325 186.680 676.000 190.720 ;
        RECT 14.325 185.280 675.600 186.680 ;
        RECT 14.325 181.920 676.000 185.280 ;
        RECT 14.325 180.520 675.600 181.920 ;
        RECT 14.325 176.480 676.000 180.520 ;
        RECT 14.325 175.080 675.600 176.480 ;
        RECT 14.325 171.720 676.000 175.080 ;
        RECT 14.325 170.320 675.600 171.720 ;
        RECT 14.325 166.280 676.000 170.320 ;
        RECT 14.325 164.880 675.600 166.280 ;
        RECT 14.325 161.520 676.000 164.880 ;
        RECT 14.325 160.120 675.600 161.520 ;
        RECT 14.325 156.080 676.000 160.120 ;
        RECT 14.325 154.680 675.600 156.080 ;
        RECT 14.325 151.320 676.000 154.680 ;
        RECT 14.325 149.920 675.600 151.320 ;
        RECT 14.325 145.880 676.000 149.920 ;
        RECT 14.325 144.480 675.600 145.880 ;
        RECT 14.325 141.120 676.000 144.480 ;
        RECT 14.325 139.720 675.600 141.120 ;
        RECT 14.325 135.680 676.000 139.720 ;
        RECT 14.325 134.280 675.600 135.680 ;
        RECT 14.325 130.240 676.000 134.280 ;
        RECT 14.325 128.840 675.600 130.240 ;
        RECT 14.325 125.480 676.000 128.840 ;
        RECT 14.325 124.080 675.600 125.480 ;
        RECT 14.325 120.040 676.000 124.080 ;
        RECT 14.325 118.640 675.600 120.040 ;
        RECT 14.325 115.280 676.000 118.640 ;
        RECT 14.325 113.880 675.600 115.280 ;
        RECT 14.325 109.840 676.000 113.880 ;
        RECT 14.325 108.440 675.600 109.840 ;
        RECT 14.325 105.080 676.000 108.440 ;
        RECT 14.325 103.680 675.600 105.080 ;
        RECT 14.325 99.640 676.000 103.680 ;
        RECT 14.325 98.240 675.600 99.640 ;
        RECT 14.325 94.880 676.000 98.240 ;
        RECT 14.325 93.480 675.600 94.880 ;
        RECT 14.325 89.440 676.000 93.480 ;
        RECT 14.325 88.040 675.600 89.440 ;
        RECT 14.325 84.680 676.000 88.040 ;
        RECT 14.325 83.280 675.600 84.680 ;
        RECT 14.325 79.240 676.000 83.280 ;
        RECT 14.325 77.840 675.600 79.240 ;
        RECT 14.325 74.480 676.000 77.840 ;
        RECT 14.325 73.080 675.600 74.480 ;
        RECT 14.325 69.040 676.000 73.080 ;
        RECT 14.325 67.640 675.600 69.040 ;
        RECT 14.325 64.280 676.000 67.640 ;
        RECT 14.325 62.880 675.600 64.280 ;
        RECT 14.325 58.840 676.000 62.880 ;
        RECT 14.325 57.440 675.600 58.840 ;
        RECT 14.325 54.080 676.000 57.440 ;
        RECT 14.325 52.680 675.600 54.080 ;
        RECT 14.325 48.640 676.000 52.680 ;
        RECT 14.325 47.240 675.600 48.640 ;
        RECT 14.325 43.880 676.000 47.240 ;
        RECT 14.325 42.480 675.600 43.880 ;
        RECT 14.325 38.440 676.000 42.480 ;
        RECT 14.325 37.040 675.600 38.440 ;
        RECT 14.325 33.680 676.000 37.040 ;
        RECT 14.325 32.280 675.600 33.680 ;
        RECT 14.325 28.240 676.000 32.280 ;
        RECT 14.325 26.840 675.600 28.240 ;
        RECT 14.325 23.480 676.000 26.840 ;
        RECT 14.325 22.080 675.600 23.480 ;
        RECT 14.325 18.040 676.000 22.080 ;
        RECT 14.325 16.640 675.600 18.040 ;
        RECT 14.325 13.280 676.000 16.640 ;
        RECT 14.325 11.880 675.600 13.280 ;
        RECT 14.325 7.840 676.000 11.880 ;
        RECT 14.325 6.440 675.600 7.840 ;
        RECT 14.325 3.080 676.000 6.440 ;
        RECT 14.325 2.215 675.600 3.080 ;
      LAYER met4 ;
        RECT 34.335 17.175 97.440 664.865 ;
        RECT 99.840 17.175 174.240 664.865 ;
        RECT 176.640 17.175 251.040 664.865 ;
        RECT 253.440 17.175 327.840 664.865 ;
        RECT 330.240 17.175 404.640 664.865 ;
        RECT 407.040 17.175 481.440 664.865 ;
        RECT 483.840 17.175 558.240 664.865 ;
        RECT 560.640 17.175 635.040 664.865 ;
        RECT 637.440 17.175 662.105 664.865 ;
  END
END icache
END LIBRARY

