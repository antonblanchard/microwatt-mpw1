magic
tech sky130A
magscale 1 2
timestamp 1612121563
<< obsli1 >>
rect 1104 1377 134872 133841
<< obsm1 >>
rect 382 8 135594 133952
<< metal2 >>
rect 386 135200 442 136000
rect 1122 135200 1178 136000
rect 1950 135200 2006 136000
rect 2686 135200 2742 136000
rect 3514 135200 3570 136000
rect 4250 135200 4306 136000
rect 5078 135200 5134 136000
rect 5814 135200 5870 136000
rect 6642 135200 6698 136000
rect 7378 135200 7434 136000
rect 8206 135200 8262 136000
rect 8942 135200 8998 136000
rect 9770 135200 9826 136000
rect 10598 135200 10654 136000
rect 11334 135200 11390 136000
rect 12162 135200 12218 136000
rect 12898 135200 12954 136000
rect 13726 135200 13782 136000
rect 14462 135200 14518 136000
rect 15290 135200 15346 136000
rect 16026 135200 16082 136000
rect 16854 135200 16910 136000
rect 17590 135200 17646 136000
rect 18418 135200 18474 136000
rect 19246 135200 19302 136000
rect 19982 135200 20038 136000
rect 20810 135200 20866 136000
rect 21546 135200 21602 136000
rect 22374 135200 22430 136000
rect 23110 135200 23166 136000
rect 23938 135200 23994 136000
rect 24674 135200 24730 136000
rect 25502 135200 25558 136000
rect 26238 135200 26294 136000
rect 27066 135200 27122 136000
rect 27894 135200 27950 136000
rect 28630 135200 28686 136000
rect 29458 135200 29514 136000
rect 30194 135200 30250 136000
rect 31022 135200 31078 136000
rect 31758 135200 31814 136000
rect 32586 135200 32642 136000
rect 33322 135200 33378 136000
rect 34150 135200 34206 136000
rect 34886 135200 34942 136000
rect 35714 135200 35770 136000
rect 36450 135200 36506 136000
rect 37278 135200 37334 136000
rect 38106 135200 38162 136000
rect 38842 135200 38898 136000
rect 39670 135200 39726 136000
rect 40406 135200 40462 136000
rect 41234 135200 41290 136000
rect 41970 135200 42026 136000
rect 42798 135200 42854 136000
rect 43534 135200 43590 136000
rect 44362 135200 44418 136000
rect 45098 135200 45154 136000
rect 45926 135200 45982 136000
rect 46754 135200 46810 136000
rect 47490 135200 47546 136000
rect 48318 135200 48374 136000
rect 49054 135200 49110 136000
rect 49882 135200 49938 136000
rect 50618 135200 50674 136000
rect 51446 135200 51502 136000
rect 52182 135200 52238 136000
rect 53010 135200 53066 136000
rect 53746 135200 53802 136000
rect 54574 135200 54630 136000
rect 55402 135200 55458 136000
rect 56138 135200 56194 136000
rect 56966 135200 57022 136000
rect 57702 135200 57758 136000
rect 58530 135200 58586 136000
rect 59266 135200 59322 136000
rect 60094 135200 60150 136000
rect 60830 135200 60886 136000
rect 61658 135200 61714 136000
rect 62394 135200 62450 136000
rect 63222 135200 63278 136000
rect 64050 135200 64106 136000
rect 64786 135200 64842 136000
rect 65614 135200 65670 136000
rect 66350 135200 66406 136000
rect 67178 135200 67234 136000
rect 67914 135200 67970 136000
rect 68742 135200 68798 136000
rect 69478 135200 69534 136000
rect 70306 135200 70362 136000
rect 71042 135200 71098 136000
rect 71870 135200 71926 136000
rect 72606 135200 72662 136000
rect 73434 135200 73490 136000
rect 74262 135200 74318 136000
rect 74998 135200 75054 136000
rect 75826 135200 75882 136000
rect 76562 135200 76618 136000
rect 77390 135200 77446 136000
rect 78126 135200 78182 136000
rect 78954 135200 79010 136000
rect 79690 135200 79746 136000
rect 80518 135200 80574 136000
rect 81254 135200 81310 136000
rect 82082 135200 82138 136000
rect 82910 135200 82966 136000
rect 83646 135200 83702 136000
rect 84474 135200 84530 136000
rect 85210 135200 85266 136000
rect 86038 135200 86094 136000
rect 86774 135200 86830 136000
rect 87602 135200 87658 136000
rect 88338 135200 88394 136000
rect 89166 135200 89222 136000
rect 89902 135200 89958 136000
rect 90730 135200 90786 136000
rect 91558 135200 91614 136000
rect 92294 135200 92350 136000
rect 93122 135200 93178 136000
rect 93858 135200 93914 136000
rect 94686 135200 94742 136000
rect 95422 135200 95478 136000
rect 96250 135200 96306 136000
rect 96986 135200 97042 136000
rect 97814 135200 97870 136000
rect 98550 135200 98606 136000
rect 99378 135200 99434 136000
rect 100206 135200 100262 136000
rect 100942 135200 100998 136000
rect 101770 135200 101826 136000
rect 102506 135200 102562 136000
rect 103334 135200 103390 136000
rect 104070 135200 104126 136000
rect 104898 135200 104954 136000
rect 105634 135200 105690 136000
rect 106462 135200 106518 136000
rect 107198 135200 107254 136000
rect 108026 135200 108082 136000
rect 108762 135200 108818 136000
rect 109590 135200 109646 136000
rect 110418 135200 110474 136000
rect 111154 135200 111210 136000
rect 111982 135200 112038 136000
rect 112718 135200 112774 136000
rect 113546 135200 113602 136000
rect 114282 135200 114338 136000
rect 115110 135200 115166 136000
rect 115846 135200 115902 136000
rect 116674 135200 116730 136000
rect 117410 135200 117466 136000
rect 118238 135200 118294 136000
rect 119066 135200 119122 136000
rect 119802 135200 119858 136000
rect 120630 135200 120686 136000
rect 121366 135200 121422 136000
rect 122194 135200 122250 136000
rect 122930 135200 122986 136000
rect 123758 135200 123814 136000
rect 124494 135200 124550 136000
rect 125322 135200 125378 136000
rect 126058 135200 126114 136000
rect 126886 135200 126942 136000
rect 127714 135200 127770 136000
rect 128450 135200 128506 136000
rect 129278 135200 129334 136000
rect 130014 135200 130070 136000
rect 130842 135200 130898 136000
rect 131578 135200 131634 136000
rect 132406 135200 132462 136000
rect 133142 135200 133198 136000
rect 133970 135200 134026 136000
rect 134706 135200 134762 136000
rect 135534 135200 135590 136000
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2686 0 2742 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 5078 0 5134 800
rect 5814 0 5870 800
rect 6642 0 6698 800
rect 7378 0 7434 800
rect 8206 0 8262 800
rect 8942 0 8998 800
rect 9770 0 9826 800
rect 10598 0 10654 800
rect 11334 0 11390 800
rect 12162 0 12218 800
rect 12898 0 12954 800
rect 13726 0 13782 800
rect 14462 0 14518 800
rect 15290 0 15346 800
rect 16026 0 16082 800
rect 16854 0 16910 800
rect 17590 0 17646 800
rect 18418 0 18474 800
rect 19246 0 19302 800
rect 19982 0 20038 800
rect 20810 0 20866 800
rect 21546 0 21602 800
rect 22374 0 22430 800
rect 23110 0 23166 800
rect 23938 0 23994 800
rect 24674 0 24730 800
rect 25502 0 25558 800
rect 26238 0 26294 800
rect 27066 0 27122 800
rect 27894 0 27950 800
rect 28630 0 28686 800
rect 29458 0 29514 800
rect 30194 0 30250 800
rect 31022 0 31078 800
rect 31758 0 31814 800
rect 32586 0 32642 800
rect 33322 0 33378 800
rect 34150 0 34206 800
rect 34886 0 34942 800
rect 35714 0 35770 800
rect 36450 0 36506 800
rect 37278 0 37334 800
rect 38106 0 38162 800
rect 38842 0 38898 800
rect 39670 0 39726 800
rect 40406 0 40462 800
rect 41234 0 41290 800
rect 41970 0 42026 800
rect 42798 0 42854 800
rect 43534 0 43590 800
rect 44362 0 44418 800
rect 45098 0 45154 800
rect 45926 0 45982 800
rect 46754 0 46810 800
rect 47490 0 47546 800
rect 48318 0 48374 800
rect 49054 0 49110 800
rect 49882 0 49938 800
rect 50618 0 50674 800
rect 51446 0 51502 800
rect 52182 0 52238 800
rect 53010 0 53066 800
rect 53746 0 53802 800
rect 54574 0 54630 800
rect 55402 0 55458 800
rect 56138 0 56194 800
rect 56966 0 57022 800
rect 57702 0 57758 800
rect 58530 0 58586 800
rect 59266 0 59322 800
rect 60094 0 60150 800
rect 60830 0 60886 800
rect 61658 0 61714 800
rect 62394 0 62450 800
rect 63222 0 63278 800
rect 64050 0 64106 800
rect 64786 0 64842 800
rect 65614 0 65670 800
rect 66350 0 66406 800
rect 67178 0 67234 800
rect 67914 0 67970 800
rect 68742 0 68798 800
rect 69478 0 69534 800
rect 70306 0 70362 800
rect 71042 0 71098 800
rect 71870 0 71926 800
rect 72606 0 72662 800
rect 73434 0 73490 800
rect 74262 0 74318 800
rect 74998 0 75054 800
rect 75826 0 75882 800
rect 76562 0 76618 800
rect 77390 0 77446 800
rect 78126 0 78182 800
rect 78954 0 79010 800
rect 79690 0 79746 800
rect 80518 0 80574 800
rect 81254 0 81310 800
rect 82082 0 82138 800
rect 82910 0 82966 800
rect 83646 0 83702 800
rect 84474 0 84530 800
rect 85210 0 85266 800
rect 86038 0 86094 800
rect 86774 0 86830 800
rect 87602 0 87658 800
rect 88338 0 88394 800
rect 89166 0 89222 800
rect 89902 0 89958 800
rect 90730 0 90786 800
rect 91558 0 91614 800
rect 92294 0 92350 800
rect 93122 0 93178 800
rect 93858 0 93914 800
rect 94686 0 94742 800
rect 95422 0 95478 800
rect 96250 0 96306 800
rect 96986 0 97042 800
rect 97814 0 97870 800
rect 98550 0 98606 800
rect 99378 0 99434 800
rect 100206 0 100262 800
rect 100942 0 100998 800
rect 101770 0 101826 800
rect 102506 0 102562 800
rect 103334 0 103390 800
rect 104070 0 104126 800
rect 104898 0 104954 800
rect 105634 0 105690 800
rect 106462 0 106518 800
rect 107198 0 107254 800
rect 108026 0 108082 800
rect 108762 0 108818 800
rect 109590 0 109646 800
rect 110418 0 110474 800
rect 111154 0 111210 800
rect 111982 0 112038 800
rect 112718 0 112774 800
rect 113546 0 113602 800
rect 114282 0 114338 800
rect 115110 0 115166 800
rect 115846 0 115902 800
rect 116674 0 116730 800
rect 117410 0 117466 800
rect 118238 0 118294 800
rect 119066 0 119122 800
rect 119802 0 119858 800
rect 120630 0 120686 800
rect 121366 0 121422 800
rect 122194 0 122250 800
rect 122930 0 122986 800
rect 123758 0 123814 800
rect 124494 0 124550 800
rect 125322 0 125378 800
rect 126058 0 126114 800
rect 126886 0 126942 800
rect 127714 0 127770 800
rect 128450 0 128506 800
rect 129278 0 129334 800
rect 130014 0 130070 800
rect 130842 0 130898 800
rect 131578 0 131634 800
rect 132406 0 132462 800
rect 133142 0 133198 800
rect 133970 0 134026 800
rect 134706 0 134762 800
rect 135534 0 135590 800
<< obsm2 >>
rect 498 135144 1066 135200
rect 1234 135144 1894 135200
rect 2062 135144 2630 135200
rect 2798 135144 3458 135200
rect 3626 135144 4194 135200
rect 4362 135144 5022 135200
rect 5190 135144 5758 135200
rect 5926 135144 6586 135200
rect 6754 135144 7322 135200
rect 7490 135144 8150 135200
rect 8318 135144 8886 135200
rect 9054 135144 9714 135200
rect 9882 135144 10542 135200
rect 10710 135144 11278 135200
rect 11446 135144 12106 135200
rect 12274 135144 12842 135200
rect 13010 135144 13670 135200
rect 13838 135144 14406 135200
rect 14574 135144 15234 135200
rect 15402 135144 15970 135200
rect 16138 135144 16798 135200
rect 16966 135144 17534 135200
rect 17702 135144 18362 135200
rect 18530 135144 19190 135200
rect 19358 135144 19926 135200
rect 20094 135144 20754 135200
rect 20922 135144 21490 135200
rect 21658 135144 22318 135200
rect 22486 135144 23054 135200
rect 23222 135144 23882 135200
rect 24050 135144 24618 135200
rect 24786 135144 25446 135200
rect 25614 135144 26182 135200
rect 26350 135144 27010 135200
rect 27178 135144 27838 135200
rect 28006 135144 28574 135200
rect 28742 135144 29402 135200
rect 29570 135144 30138 135200
rect 30306 135144 30966 135200
rect 31134 135144 31702 135200
rect 31870 135144 32530 135200
rect 32698 135144 33266 135200
rect 33434 135144 34094 135200
rect 34262 135144 34830 135200
rect 34998 135144 35658 135200
rect 35826 135144 36394 135200
rect 36562 135144 37222 135200
rect 37390 135144 38050 135200
rect 38218 135144 38786 135200
rect 38954 135144 39614 135200
rect 39782 135144 40350 135200
rect 40518 135144 41178 135200
rect 41346 135144 41914 135200
rect 42082 135144 42742 135200
rect 42910 135144 43478 135200
rect 43646 135144 44306 135200
rect 44474 135144 45042 135200
rect 45210 135144 45870 135200
rect 46038 135144 46698 135200
rect 46866 135144 47434 135200
rect 47602 135144 48262 135200
rect 48430 135144 48998 135200
rect 49166 135144 49826 135200
rect 49994 135144 50562 135200
rect 50730 135144 51390 135200
rect 51558 135144 52126 135200
rect 52294 135144 52954 135200
rect 53122 135144 53690 135200
rect 53858 135144 54518 135200
rect 54686 135144 55346 135200
rect 55514 135144 56082 135200
rect 56250 135144 56910 135200
rect 57078 135144 57646 135200
rect 57814 135144 58474 135200
rect 58642 135144 59210 135200
rect 59378 135144 60038 135200
rect 60206 135144 60774 135200
rect 60942 135144 61602 135200
rect 61770 135144 62338 135200
rect 62506 135144 63166 135200
rect 63334 135144 63994 135200
rect 64162 135144 64730 135200
rect 64898 135144 65558 135200
rect 65726 135144 66294 135200
rect 66462 135144 67122 135200
rect 67290 135144 67858 135200
rect 68026 135144 68686 135200
rect 68854 135144 69422 135200
rect 69590 135144 70250 135200
rect 70418 135144 70986 135200
rect 71154 135144 71814 135200
rect 71982 135144 72550 135200
rect 72718 135144 73378 135200
rect 73546 135144 74206 135200
rect 74374 135144 74942 135200
rect 75110 135144 75770 135200
rect 75938 135144 76506 135200
rect 76674 135144 77334 135200
rect 77502 135144 78070 135200
rect 78238 135144 78898 135200
rect 79066 135144 79634 135200
rect 79802 135144 80462 135200
rect 80630 135144 81198 135200
rect 81366 135144 82026 135200
rect 82194 135144 82854 135200
rect 83022 135144 83590 135200
rect 83758 135144 84418 135200
rect 84586 135144 85154 135200
rect 85322 135144 85982 135200
rect 86150 135144 86718 135200
rect 86886 135144 87546 135200
rect 87714 135144 88282 135200
rect 88450 135144 89110 135200
rect 89278 135144 89846 135200
rect 90014 135144 90674 135200
rect 90842 135144 91502 135200
rect 91670 135144 92238 135200
rect 92406 135144 93066 135200
rect 93234 135144 93802 135200
rect 93970 135144 94630 135200
rect 94798 135144 95366 135200
rect 95534 135144 96194 135200
rect 96362 135144 96930 135200
rect 97098 135144 97758 135200
rect 97926 135144 98494 135200
rect 98662 135144 99322 135200
rect 99490 135144 100150 135200
rect 100318 135144 100886 135200
rect 101054 135144 101714 135200
rect 101882 135144 102450 135200
rect 102618 135144 103278 135200
rect 103446 135144 104014 135200
rect 104182 135144 104842 135200
rect 105010 135144 105578 135200
rect 105746 135144 106406 135200
rect 106574 135144 107142 135200
rect 107310 135144 107970 135200
rect 108138 135144 108706 135200
rect 108874 135144 109534 135200
rect 109702 135144 110362 135200
rect 110530 135144 111098 135200
rect 111266 135144 111926 135200
rect 112094 135144 112662 135200
rect 112830 135144 113490 135200
rect 113658 135144 114226 135200
rect 114394 135144 115054 135200
rect 115222 135144 115790 135200
rect 115958 135144 116618 135200
rect 116786 135144 117354 135200
rect 117522 135144 118182 135200
rect 118350 135144 119010 135200
rect 119178 135144 119746 135200
rect 119914 135144 120574 135200
rect 120742 135144 121310 135200
rect 121478 135144 122138 135200
rect 122306 135144 122874 135200
rect 123042 135144 123702 135200
rect 123870 135144 124438 135200
rect 124606 135144 125266 135200
rect 125434 135144 126002 135200
rect 126170 135144 126830 135200
rect 126998 135144 127658 135200
rect 127826 135144 128394 135200
rect 128562 135144 129222 135200
rect 129390 135144 129958 135200
rect 130126 135144 130786 135200
rect 130954 135144 131522 135200
rect 131690 135144 132350 135200
rect 132518 135144 133086 135200
rect 133254 135144 133914 135200
rect 134082 135144 134650 135200
rect 134818 135144 135478 135200
rect 388 856 135588 135144
rect 498 2 1066 856
rect 1234 2 1894 856
rect 2062 2 2630 856
rect 2798 2 3458 856
rect 3626 2 4194 856
rect 4362 2 5022 856
rect 5190 2 5758 856
rect 5926 2 6586 856
rect 6754 2 7322 856
rect 7490 2 8150 856
rect 8318 2 8886 856
rect 9054 2 9714 856
rect 9882 2 10542 856
rect 10710 2 11278 856
rect 11446 2 12106 856
rect 12274 2 12842 856
rect 13010 2 13670 856
rect 13838 2 14406 856
rect 14574 2 15234 856
rect 15402 2 15970 856
rect 16138 2 16798 856
rect 16966 2 17534 856
rect 17702 2 18362 856
rect 18530 2 19190 856
rect 19358 2 19926 856
rect 20094 2 20754 856
rect 20922 2 21490 856
rect 21658 2 22318 856
rect 22486 2 23054 856
rect 23222 2 23882 856
rect 24050 2 24618 856
rect 24786 2 25446 856
rect 25614 2 26182 856
rect 26350 2 27010 856
rect 27178 2 27838 856
rect 28006 2 28574 856
rect 28742 2 29402 856
rect 29570 2 30138 856
rect 30306 2 30966 856
rect 31134 2 31702 856
rect 31870 2 32530 856
rect 32698 2 33266 856
rect 33434 2 34094 856
rect 34262 2 34830 856
rect 34998 2 35658 856
rect 35826 2 36394 856
rect 36562 2 37222 856
rect 37390 2 38050 856
rect 38218 2 38786 856
rect 38954 2 39614 856
rect 39782 2 40350 856
rect 40518 2 41178 856
rect 41346 2 41914 856
rect 42082 2 42742 856
rect 42910 2 43478 856
rect 43646 2 44306 856
rect 44474 2 45042 856
rect 45210 2 45870 856
rect 46038 2 46698 856
rect 46866 2 47434 856
rect 47602 2 48262 856
rect 48430 2 48998 856
rect 49166 2 49826 856
rect 49994 2 50562 856
rect 50730 2 51390 856
rect 51558 2 52126 856
rect 52294 2 52954 856
rect 53122 2 53690 856
rect 53858 2 54518 856
rect 54686 2 55346 856
rect 55514 2 56082 856
rect 56250 2 56910 856
rect 57078 2 57646 856
rect 57814 2 58474 856
rect 58642 2 59210 856
rect 59378 2 60038 856
rect 60206 2 60774 856
rect 60942 2 61602 856
rect 61770 2 62338 856
rect 62506 2 63166 856
rect 63334 2 63994 856
rect 64162 2 64730 856
rect 64898 2 65558 856
rect 65726 2 66294 856
rect 66462 2 67122 856
rect 67290 2 67858 856
rect 68026 2 68686 856
rect 68854 2 69422 856
rect 69590 2 70250 856
rect 70418 2 70986 856
rect 71154 2 71814 856
rect 71982 2 72550 856
rect 72718 2 73378 856
rect 73546 2 74206 856
rect 74374 2 74942 856
rect 75110 2 75770 856
rect 75938 2 76506 856
rect 76674 2 77334 856
rect 77502 2 78070 856
rect 78238 2 78898 856
rect 79066 2 79634 856
rect 79802 2 80462 856
rect 80630 2 81198 856
rect 81366 2 82026 856
rect 82194 2 82854 856
rect 83022 2 83590 856
rect 83758 2 84418 856
rect 84586 2 85154 856
rect 85322 2 85982 856
rect 86150 2 86718 856
rect 86886 2 87546 856
rect 87714 2 88282 856
rect 88450 2 89110 856
rect 89278 2 89846 856
rect 90014 2 90674 856
rect 90842 2 91502 856
rect 91670 2 92238 856
rect 92406 2 93066 856
rect 93234 2 93802 856
rect 93970 2 94630 856
rect 94798 2 95366 856
rect 95534 2 96194 856
rect 96362 2 96930 856
rect 97098 2 97758 856
rect 97926 2 98494 856
rect 98662 2 99322 856
rect 99490 2 100150 856
rect 100318 2 100886 856
rect 101054 2 101714 856
rect 101882 2 102450 856
rect 102618 2 103278 856
rect 103446 2 104014 856
rect 104182 2 104842 856
rect 105010 2 105578 856
rect 105746 2 106406 856
rect 106574 2 107142 856
rect 107310 2 107970 856
rect 108138 2 108706 856
rect 108874 2 109534 856
rect 109702 2 110362 856
rect 110530 2 111098 856
rect 111266 2 111926 856
rect 112094 2 112662 856
rect 112830 2 113490 856
rect 113658 2 114226 856
rect 114394 2 115054 856
rect 115222 2 115790 856
rect 115958 2 116618 856
rect 116786 2 117354 856
rect 117522 2 118182 856
rect 118350 2 119010 856
rect 119178 2 119746 856
rect 119914 2 120574 856
rect 120742 2 121310 856
rect 121478 2 122138 856
rect 122306 2 122874 856
rect 123042 2 123702 856
rect 123870 2 124438 856
rect 124606 2 125266 856
rect 125434 2 126002 856
rect 126170 2 126830 856
rect 126998 2 127658 856
rect 127826 2 128394 856
rect 128562 2 129222 856
rect 129390 2 129958 856
rect 130126 2 130786 856
rect 130954 2 131522 856
rect 131690 2 132350 856
rect 132518 2 133086 856
rect 133254 2 133914 856
rect 134082 2 134650 856
rect 134818 2 135478 856
<< metal3 >>
rect 135200 135328 136000 135448
rect 135200 134240 136000 134360
rect 135200 133288 136000 133408
rect 135200 132200 136000 132320
rect 135200 131248 136000 131368
rect 135200 130160 136000 130280
rect 135200 129208 136000 129328
rect 135200 128120 136000 128240
rect 135200 127168 136000 127288
rect 135200 126080 136000 126200
rect 135200 125128 136000 125248
rect 135200 124040 136000 124160
rect 135200 123088 136000 123208
rect 135200 122000 136000 122120
rect 135200 121048 136000 121168
rect 135200 119960 136000 120080
rect 135200 119008 136000 119128
rect 135200 117920 136000 118040
rect 135200 116968 136000 117088
rect 135200 115880 136000 116000
rect 135200 114928 136000 115048
rect 135200 113840 136000 113960
rect 135200 112888 136000 113008
rect 135200 111800 136000 111920
rect 135200 110848 136000 110968
rect 135200 109760 136000 109880
rect 135200 108672 136000 108792
rect 135200 107720 136000 107840
rect 135200 106632 136000 106752
rect 135200 105680 136000 105800
rect 135200 104592 136000 104712
rect 135200 103640 136000 103760
rect 135200 102552 136000 102672
rect 135200 101600 136000 101720
rect 135200 100512 136000 100632
rect 135200 99560 136000 99680
rect 135200 98472 136000 98592
rect 135200 97520 136000 97640
rect 135200 96432 136000 96552
rect 135200 95480 136000 95600
rect 135200 94392 136000 94512
rect 135200 93440 136000 93560
rect 135200 92352 136000 92472
rect 135200 91400 136000 91520
rect 135200 90312 136000 90432
rect 135200 89360 136000 89480
rect 135200 88272 136000 88392
rect 135200 87320 136000 87440
rect 135200 86232 136000 86352
rect 135200 85280 136000 85400
rect 135200 84192 136000 84312
rect 135200 83240 136000 83360
rect 135200 82152 136000 82272
rect 135200 81064 136000 81184
rect 135200 80112 136000 80232
rect 135200 79024 136000 79144
rect 135200 78072 136000 78192
rect 135200 76984 136000 77104
rect 135200 76032 136000 76152
rect 135200 74944 136000 75064
rect 135200 73992 136000 74112
rect 135200 72904 136000 73024
rect 135200 71952 136000 72072
rect 135200 70864 136000 70984
rect 135200 69912 136000 70032
rect 135200 68824 136000 68944
rect 135200 67872 136000 67992
rect 135200 66784 136000 66904
rect 135200 65832 136000 65952
rect 135200 64744 136000 64864
rect 135200 63792 136000 63912
rect 135200 62704 136000 62824
rect 135200 61752 136000 61872
rect 135200 60664 136000 60784
rect 135200 59712 136000 59832
rect 135200 58624 136000 58744
rect 135200 57672 136000 57792
rect 135200 56584 136000 56704
rect 135200 55632 136000 55752
rect 135200 54544 136000 54664
rect 135200 53456 136000 53576
rect 135200 52504 136000 52624
rect 135200 51416 136000 51536
rect 135200 50464 136000 50584
rect 135200 49376 136000 49496
rect 135200 48424 136000 48544
rect 135200 47336 136000 47456
rect 135200 46384 136000 46504
rect 135200 45296 136000 45416
rect 135200 44344 136000 44464
rect 135200 43256 136000 43376
rect 135200 42304 136000 42424
rect 135200 41216 136000 41336
rect 135200 40264 136000 40384
rect 135200 39176 136000 39296
rect 135200 38224 136000 38344
rect 135200 37136 136000 37256
rect 135200 36184 136000 36304
rect 135200 35096 136000 35216
rect 135200 34144 136000 34264
rect 135200 33056 136000 33176
rect 135200 32104 136000 32224
rect 135200 31016 136000 31136
rect 135200 30064 136000 30184
rect 135200 28976 136000 29096
rect 135200 28024 136000 28144
rect 135200 26936 136000 27056
rect 135200 25848 136000 25968
rect 135200 24896 136000 25016
rect 135200 23808 136000 23928
rect 135200 22856 136000 22976
rect 135200 21768 136000 21888
rect 135200 20816 136000 20936
rect 135200 19728 136000 19848
rect 135200 18776 136000 18896
rect 135200 17688 136000 17808
rect 135200 16736 136000 16856
rect 135200 15648 136000 15768
rect 135200 14696 136000 14816
rect 135200 13608 136000 13728
rect 135200 12656 136000 12776
rect 135200 11568 136000 11688
rect 135200 10616 136000 10736
rect 135200 9528 136000 9648
rect 135200 8576 136000 8696
rect 135200 7488 136000 7608
rect 135200 6536 136000 6656
rect 135200 5448 136000 5568
rect 135200 4496 136000 4616
rect 135200 3408 136000 3528
rect 135200 2456 136000 2576
rect 135200 1368 136000 1488
rect 135200 416 136000 536
<< obsm3 >>
rect 2865 133488 135200 133857
rect 2865 133208 135120 133488
rect 2865 132400 135200 133208
rect 2865 132120 135120 132400
rect 2865 131448 135200 132120
rect 2865 131168 135120 131448
rect 2865 130360 135200 131168
rect 2865 130080 135120 130360
rect 2865 129408 135200 130080
rect 2865 129128 135120 129408
rect 2865 128320 135200 129128
rect 2865 128040 135120 128320
rect 2865 127368 135200 128040
rect 2865 127088 135120 127368
rect 2865 126280 135200 127088
rect 2865 126000 135120 126280
rect 2865 125328 135200 126000
rect 2865 125048 135120 125328
rect 2865 124240 135200 125048
rect 2865 123960 135120 124240
rect 2865 123288 135200 123960
rect 2865 123008 135120 123288
rect 2865 122200 135200 123008
rect 2865 121920 135120 122200
rect 2865 121248 135200 121920
rect 2865 120968 135120 121248
rect 2865 120160 135200 120968
rect 2865 119880 135120 120160
rect 2865 119208 135200 119880
rect 2865 118928 135120 119208
rect 2865 118120 135200 118928
rect 2865 117840 135120 118120
rect 2865 117168 135200 117840
rect 2865 116888 135120 117168
rect 2865 116080 135200 116888
rect 2865 115800 135120 116080
rect 2865 115128 135200 115800
rect 2865 114848 135120 115128
rect 2865 114040 135200 114848
rect 2865 113760 135120 114040
rect 2865 113088 135200 113760
rect 2865 112808 135120 113088
rect 2865 112000 135200 112808
rect 2865 111720 135120 112000
rect 2865 111048 135200 111720
rect 2865 110768 135120 111048
rect 2865 109960 135200 110768
rect 2865 109680 135120 109960
rect 2865 108872 135200 109680
rect 2865 108592 135120 108872
rect 2865 107920 135200 108592
rect 2865 107640 135120 107920
rect 2865 106832 135200 107640
rect 2865 106552 135120 106832
rect 2865 105880 135200 106552
rect 2865 105600 135120 105880
rect 2865 104792 135200 105600
rect 2865 104512 135120 104792
rect 2865 103840 135200 104512
rect 2865 103560 135120 103840
rect 2865 102752 135200 103560
rect 2865 102472 135120 102752
rect 2865 101800 135200 102472
rect 2865 101520 135120 101800
rect 2865 100712 135200 101520
rect 2865 100432 135120 100712
rect 2865 99760 135200 100432
rect 2865 99480 135120 99760
rect 2865 98672 135200 99480
rect 2865 98392 135120 98672
rect 2865 97720 135200 98392
rect 2865 97440 135120 97720
rect 2865 96632 135200 97440
rect 2865 96352 135120 96632
rect 2865 95680 135200 96352
rect 2865 95400 135120 95680
rect 2865 94592 135200 95400
rect 2865 94312 135120 94592
rect 2865 93640 135200 94312
rect 2865 93360 135120 93640
rect 2865 92552 135200 93360
rect 2865 92272 135120 92552
rect 2865 91600 135200 92272
rect 2865 91320 135120 91600
rect 2865 90512 135200 91320
rect 2865 90232 135120 90512
rect 2865 89560 135200 90232
rect 2865 89280 135120 89560
rect 2865 88472 135200 89280
rect 2865 88192 135120 88472
rect 2865 87520 135200 88192
rect 2865 87240 135120 87520
rect 2865 86432 135200 87240
rect 2865 86152 135120 86432
rect 2865 85480 135200 86152
rect 2865 85200 135120 85480
rect 2865 84392 135200 85200
rect 2865 84112 135120 84392
rect 2865 83440 135200 84112
rect 2865 83160 135120 83440
rect 2865 82352 135200 83160
rect 2865 82072 135120 82352
rect 2865 81264 135200 82072
rect 2865 80984 135120 81264
rect 2865 80312 135200 80984
rect 2865 80032 135120 80312
rect 2865 79224 135200 80032
rect 2865 78944 135120 79224
rect 2865 78272 135200 78944
rect 2865 77992 135120 78272
rect 2865 77184 135200 77992
rect 2865 76904 135120 77184
rect 2865 76232 135200 76904
rect 2865 75952 135120 76232
rect 2865 75144 135200 75952
rect 2865 74864 135120 75144
rect 2865 74192 135200 74864
rect 2865 73912 135120 74192
rect 2865 73104 135200 73912
rect 2865 72824 135120 73104
rect 2865 72152 135200 72824
rect 2865 71872 135120 72152
rect 2865 71064 135200 71872
rect 2865 70784 135120 71064
rect 2865 70112 135200 70784
rect 2865 69832 135120 70112
rect 2865 69024 135200 69832
rect 2865 68744 135120 69024
rect 2865 68072 135200 68744
rect 2865 67792 135120 68072
rect 2865 66984 135200 67792
rect 2865 66704 135120 66984
rect 2865 66032 135200 66704
rect 2865 65752 135120 66032
rect 2865 64944 135200 65752
rect 2865 64664 135120 64944
rect 2865 63992 135200 64664
rect 2865 63712 135120 63992
rect 2865 62904 135200 63712
rect 2865 62624 135120 62904
rect 2865 61952 135200 62624
rect 2865 61672 135120 61952
rect 2865 60864 135200 61672
rect 2865 60584 135120 60864
rect 2865 59912 135200 60584
rect 2865 59632 135120 59912
rect 2865 58824 135200 59632
rect 2865 58544 135120 58824
rect 2865 57872 135200 58544
rect 2865 57592 135120 57872
rect 2865 56784 135200 57592
rect 2865 56504 135120 56784
rect 2865 55832 135200 56504
rect 2865 55552 135120 55832
rect 2865 54744 135200 55552
rect 2865 54464 135120 54744
rect 2865 53656 135200 54464
rect 2865 53376 135120 53656
rect 2865 52704 135200 53376
rect 2865 52424 135120 52704
rect 2865 51616 135200 52424
rect 2865 51336 135120 51616
rect 2865 50664 135200 51336
rect 2865 50384 135120 50664
rect 2865 49576 135200 50384
rect 2865 49296 135120 49576
rect 2865 48624 135200 49296
rect 2865 48344 135120 48624
rect 2865 47536 135200 48344
rect 2865 47256 135120 47536
rect 2865 46584 135200 47256
rect 2865 46304 135120 46584
rect 2865 45496 135200 46304
rect 2865 45216 135120 45496
rect 2865 44544 135200 45216
rect 2865 44264 135120 44544
rect 2865 43456 135200 44264
rect 2865 43176 135120 43456
rect 2865 42504 135200 43176
rect 2865 42224 135120 42504
rect 2865 41416 135200 42224
rect 2865 41136 135120 41416
rect 2865 40464 135200 41136
rect 2865 40184 135120 40464
rect 2865 39376 135200 40184
rect 2865 39096 135120 39376
rect 2865 38424 135200 39096
rect 2865 38144 135120 38424
rect 2865 37336 135200 38144
rect 2865 37056 135120 37336
rect 2865 36384 135200 37056
rect 2865 36104 135120 36384
rect 2865 35296 135200 36104
rect 2865 35016 135120 35296
rect 2865 34344 135200 35016
rect 2865 34064 135120 34344
rect 2865 33256 135200 34064
rect 2865 32976 135120 33256
rect 2865 32304 135200 32976
rect 2865 32024 135120 32304
rect 2865 31216 135200 32024
rect 2865 30936 135120 31216
rect 2865 30264 135200 30936
rect 2865 29984 135120 30264
rect 2865 29176 135200 29984
rect 2865 28896 135120 29176
rect 2865 28224 135200 28896
rect 2865 27944 135120 28224
rect 2865 27136 135200 27944
rect 2865 26856 135120 27136
rect 2865 26048 135200 26856
rect 2865 25768 135120 26048
rect 2865 25096 135200 25768
rect 2865 24816 135120 25096
rect 2865 24008 135200 24816
rect 2865 23728 135120 24008
rect 2865 23056 135200 23728
rect 2865 22776 135120 23056
rect 2865 21968 135200 22776
rect 2865 21688 135120 21968
rect 2865 21016 135200 21688
rect 2865 20736 135120 21016
rect 2865 19928 135200 20736
rect 2865 19648 135120 19928
rect 2865 18976 135200 19648
rect 2865 18696 135120 18976
rect 2865 17888 135200 18696
rect 2865 17608 135120 17888
rect 2865 16936 135200 17608
rect 2865 16656 135120 16936
rect 2865 15848 135200 16656
rect 2865 15568 135120 15848
rect 2865 14896 135200 15568
rect 2865 14616 135120 14896
rect 2865 13808 135200 14616
rect 2865 13528 135120 13808
rect 2865 12856 135200 13528
rect 2865 12576 135120 12856
rect 2865 11768 135200 12576
rect 2865 11488 135120 11768
rect 2865 10816 135200 11488
rect 2865 10536 135120 10816
rect 2865 9728 135200 10536
rect 2865 9448 135120 9728
rect 2865 8776 135200 9448
rect 2865 8496 135120 8776
rect 2865 7688 135200 8496
rect 2865 7408 135120 7688
rect 2865 6736 135200 7408
rect 2865 6456 135120 6736
rect 2865 5648 135200 6456
rect 2865 5368 135120 5648
rect 2865 4696 135200 5368
rect 2865 4416 135120 4696
rect 2865 3608 135200 4416
rect 2865 3328 135120 3608
rect 2865 2656 135200 3328
rect 2865 2376 135120 2656
rect 2865 1568 135200 2376
rect 2865 1288 135120 1568
rect 2865 616 135200 1288
rect 2865 443 135120 616
<< metal4 >>
rect 4208 2128 4528 133872
rect 19568 2128 19888 133872
rect 34928 2128 35248 133872
rect 50288 2128 50608 133872
rect 65648 2128 65968 133872
rect 81008 2128 81328 133872
rect 96368 2128 96688 133872
rect 111728 2128 112048 133872
rect 127088 2128 127408 133872
<< obsm4 >>
rect 6867 3435 19488 132973
rect 19968 3435 34848 132973
rect 35328 3435 50208 132973
rect 50688 3435 65568 132973
rect 66048 3435 80928 132973
rect 81408 3435 96288 132973
rect 96768 3435 111648 132973
rect 112128 3435 127008 132973
rect 127488 3435 132421 132973
<< labels >>
rlabel metal3 s 135200 416 136000 536 6 clk
port 1 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 flush_in
port 2 nsew signal input
rlabel metal2 s 386 0 442 800 6 i_in[0]
port 3 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 i_in[10]
port 4 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 i_in[11]
port 5 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 i_in[12]
port 6 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 i_in[13]
port 7 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 i_in[14]
port 8 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 i_in[15]
port 9 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 i_in[16]
port 10 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 i_in[17]
port 11 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 i_in[18]
port 12 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 i_in[19]
port 13 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 i_in[1]
port 14 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 i_in[20]
port 15 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 i_in[21]
port 16 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 i_in[22]
port 17 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 i_in[23]
port 18 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 i_in[24]
port 19 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 i_in[25]
port 20 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 i_in[26]
port 21 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 i_in[27]
port 22 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 i_in[28]
port 23 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 i_in[29]
port 24 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 i_in[2]
port 25 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 i_in[30]
port 26 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 i_in[31]
port 27 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 i_in[32]
port 28 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 i_in[33]
port 29 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 i_in[34]
port 30 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 i_in[35]
port 31 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 i_in[36]
port 32 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 i_in[37]
port 33 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 i_in[38]
port 34 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 i_in[39]
port 35 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 i_in[3]
port 36 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 i_in[40]
port 37 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 i_in[41]
port 38 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 i_in[42]
port 39 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 i_in[43]
port 40 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 i_in[44]
port 41 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 i_in[45]
port 42 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 i_in[46]
port 43 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 i_in[47]
port 44 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 i_in[48]
port 45 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 i_in[49]
port 46 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 i_in[4]
port 47 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 i_in[50]
port 48 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 i_in[51]
port 49 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 i_in[52]
port 50 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 i_in[53]
port 51 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 i_in[54]
port 52 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 i_in[55]
port 53 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 i_in[56]
port 54 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 i_in[57]
port 55 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 i_in[58]
port 56 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 i_in[59]
port 57 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 i_in[5]
port 58 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 i_in[60]
port 59 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 i_in[61]
port 60 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 i_in[62]
port 61 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 i_in[63]
port 62 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 i_in[64]
port 63 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 i_in[65]
port 64 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 i_in[66]
port 65 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 i_in[67]
port 66 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 i_in[68]
port 67 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 i_in[69]
port 68 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 i_in[6]
port 69 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 i_in[7]
port 70 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 i_in[8]
port 71 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 i_in[9]
port 72 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 i_out[0]
port 73 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 i_out[10]
port 74 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 i_out[11]
port 75 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 i_out[12]
port 76 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 i_out[13]
port 77 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 i_out[14]
port 78 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 i_out[15]
port 79 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 i_out[16]
port 80 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 i_out[17]
port 81 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 i_out[18]
port 82 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 i_out[19]
port 83 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 i_out[1]
port 84 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 i_out[20]
port 85 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 i_out[21]
port 86 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 i_out[22]
port 87 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 i_out[23]
port 88 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 i_out[24]
port 89 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 i_out[25]
port 90 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 i_out[26]
port 91 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 i_out[27]
port 92 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 i_out[28]
port 93 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 i_out[29]
port 94 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 i_out[2]
port 95 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 i_out[30]
port 96 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 i_out[31]
port 97 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 i_out[32]
port 98 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 i_out[33]
port 99 nsew signal output
rlabel metal2 s 82082 0 82138 800 6 i_out[34]
port 100 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 i_out[35]
port 101 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 i_out[36]
port 102 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 i_out[37]
port 103 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 i_out[38]
port 104 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 i_out[39]
port 105 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 i_out[3]
port 106 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 i_out[40]
port 107 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 i_out[41]
port 108 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 i_out[42]
port 109 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 i_out[43]
port 110 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 i_out[44]
port 111 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 i_out[45]
port 112 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 i_out[46]
port 113 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 i_out[47]
port 114 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 i_out[48]
port 115 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 i_out[49]
port 116 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 i_out[4]
port 117 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 i_out[50]
port 118 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 i_out[51]
port 119 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 i_out[52]
port 120 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 i_out[53]
port 121 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 i_out[54]
port 122 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 i_out[55]
port 123 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 i_out[56]
port 124 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 i_out[57]
port 125 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 i_out[58]
port 126 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 i_out[59]
port 127 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 i_out[5]
port 128 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 i_out[60]
port 129 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 i_out[61]
port 130 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 i_out[62]
port 131 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 i_out[63]
port 132 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 i_out[64]
port 133 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 i_out[65]
port 134 nsew signal output
rlabel metal2 s 107198 0 107254 800 6 i_out[66]
port 135 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 i_out[67]
port 136 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 i_out[68]
port 137 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 i_out[69]
port 138 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 i_out[6]
port 139 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 i_out[70]
port 140 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 i_out[71]
port 141 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 i_out[72]
port 142 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 i_out[73]
port 143 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 i_out[74]
port 144 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 i_out[75]
port 145 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 i_out[76]
port 146 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 i_out[77]
port 147 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 i_out[78]
port 148 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 i_out[79]
port 149 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 i_out[7]
port 150 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 i_out[80]
port 151 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 i_out[81]
port 152 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 i_out[82]
port 153 nsew signal output
rlabel metal2 s 120630 0 120686 800 6 i_out[83]
port 154 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 i_out[84]
port 155 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 i_out[85]
port 156 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 i_out[86]
port 157 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 i_out[87]
port 158 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 i_out[88]
port 159 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 i_out[89]
port 160 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 i_out[8]
port 161 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 i_out[90]
port 162 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 i_out[91]
port 163 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 i_out[92]
port 164 nsew signal output
rlabel metal2 s 128450 0 128506 800 6 i_out[93]
port 165 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 i_out[94]
port 166 nsew signal output
rlabel metal2 s 130014 0 130070 800 6 i_out[95]
port 167 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 i_out[96]
port 168 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 i_out[97]
port 169 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 i_out[98]
port 170 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 i_out[9]
port 171 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 inval_in
port 172 nsew signal input
rlabel metal3 s 135200 2456 136000 2576 6 m_in[0]
port 173 nsew signal input
rlabel metal3 s 135200 104592 136000 104712 6 m_in[100]
port 174 nsew signal input
rlabel metal3 s 135200 105680 136000 105800 6 m_in[101]
port 175 nsew signal input
rlabel metal3 s 135200 106632 136000 106752 6 m_in[102]
port 176 nsew signal input
rlabel metal3 s 135200 107720 136000 107840 6 m_in[103]
port 177 nsew signal input
rlabel metal3 s 135200 108672 136000 108792 6 m_in[104]
port 178 nsew signal input
rlabel metal3 s 135200 109760 136000 109880 6 m_in[105]
port 179 nsew signal input
rlabel metal3 s 135200 110848 136000 110968 6 m_in[106]
port 180 nsew signal input
rlabel metal3 s 135200 111800 136000 111920 6 m_in[107]
port 181 nsew signal input
rlabel metal3 s 135200 112888 136000 113008 6 m_in[108]
port 182 nsew signal input
rlabel metal3 s 135200 113840 136000 113960 6 m_in[109]
port 183 nsew signal input
rlabel metal3 s 135200 12656 136000 12776 6 m_in[10]
port 184 nsew signal input
rlabel metal3 s 135200 114928 136000 115048 6 m_in[110]
port 185 nsew signal input
rlabel metal3 s 135200 115880 136000 116000 6 m_in[111]
port 186 nsew signal input
rlabel metal3 s 135200 116968 136000 117088 6 m_in[112]
port 187 nsew signal input
rlabel metal3 s 135200 117920 136000 118040 6 m_in[113]
port 188 nsew signal input
rlabel metal3 s 135200 119008 136000 119128 6 m_in[114]
port 189 nsew signal input
rlabel metal3 s 135200 119960 136000 120080 6 m_in[115]
port 190 nsew signal input
rlabel metal3 s 135200 121048 136000 121168 6 m_in[116]
port 191 nsew signal input
rlabel metal3 s 135200 122000 136000 122120 6 m_in[117]
port 192 nsew signal input
rlabel metal3 s 135200 123088 136000 123208 6 m_in[118]
port 193 nsew signal input
rlabel metal3 s 135200 124040 136000 124160 6 m_in[119]
port 194 nsew signal input
rlabel metal3 s 135200 13608 136000 13728 6 m_in[11]
port 195 nsew signal input
rlabel metal3 s 135200 125128 136000 125248 6 m_in[120]
port 196 nsew signal input
rlabel metal3 s 135200 126080 136000 126200 6 m_in[121]
port 197 nsew signal input
rlabel metal3 s 135200 127168 136000 127288 6 m_in[122]
port 198 nsew signal input
rlabel metal3 s 135200 128120 136000 128240 6 m_in[123]
port 199 nsew signal input
rlabel metal3 s 135200 129208 136000 129328 6 m_in[124]
port 200 nsew signal input
rlabel metal3 s 135200 130160 136000 130280 6 m_in[125]
port 201 nsew signal input
rlabel metal3 s 135200 131248 136000 131368 6 m_in[126]
port 202 nsew signal input
rlabel metal3 s 135200 132200 136000 132320 6 m_in[127]
port 203 nsew signal input
rlabel metal3 s 135200 133288 136000 133408 6 m_in[128]
port 204 nsew signal input
rlabel metal3 s 135200 134240 136000 134360 6 m_in[129]
port 205 nsew signal input
rlabel metal3 s 135200 14696 136000 14816 6 m_in[12]
port 206 nsew signal input
rlabel metal3 s 135200 135328 136000 135448 6 m_in[130]
port 207 nsew signal input
rlabel metal3 s 135200 15648 136000 15768 6 m_in[13]
port 208 nsew signal input
rlabel metal3 s 135200 16736 136000 16856 6 m_in[14]
port 209 nsew signal input
rlabel metal3 s 135200 17688 136000 17808 6 m_in[15]
port 210 nsew signal input
rlabel metal3 s 135200 18776 136000 18896 6 m_in[16]
port 211 nsew signal input
rlabel metal3 s 135200 19728 136000 19848 6 m_in[17]
port 212 nsew signal input
rlabel metal3 s 135200 20816 136000 20936 6 m_in[18]
port 213 nsew signal input
rlabel metal3 s 135200 21768 136000 21888 6 m_in[19]
port 214 nsew signal input
rlabel metal3 s 135200 3408 136000 3528 6 m_in[1]
port 215 nsew signal input
rlabel metal3 s 135200 22856 136000 22976 6 m_in[20]
port 216 nsew signal input
rlabel metal3 s 135200 23808 136000 23928 6 m_in[21]
port 217 nsew signal input
rlabel metal3 s 135200 24896 136000 25016 6 m_in[22]
port 218 nsew signal input
rlabel metal3 s 135200 25848 136000 25968 6 m_in[23]
port 219 nsew signal input
rlabel metal3 s 135200 26936 136000 27056 6 m_in[24]
port 220 nsew signal input
rlabel metal3 s 135200 28024 136000 28144 6 m_in[25]
port 221 nsew signal input
rlabel metal3 s 135200 28976 136000 29096 6 m_in[26]
port 222 nsew signal input
rlabel metal3 s 135200 30064 136000 30184 6 m_in[27]
port 223 nsew signal input
rlabel metal3 s 135200 31016 136000 31136 6 m_in[28]
port 224 nsew signal input
rlabel metal3 s 135200 32104 136000 32224 6 m_in[29]
port 225 nsew signal input
rlabel metal3 s 135200 4496 136000 4616 6 m_in[2]
port 226 nsew signal input
rlabel metal3 s 135200 33056 136000 33176 6 m_in[30]
port 227 nsew signal input
rlabel metal3 s 135200 34144 136000 34264 6 m_in[31]
port 228 nsew signal input
rlabel metal3 s 135200 35096 136000 35216 6 m_in[32]
port 229 nsew signal input
rlabel metal3 s 135200 36184 136000 36304 6 m_in[33]
port 230 nsew signal input
rlabel metal3 s 135200 37136 136000 37256 6 m_in[34]
port 231 nsew signal input
rlabel metal3 s 135200 38224 136000 38344 6 m_in[35]
port 232 nsew signal input
rlabel metal3 s 135200 39176 136000 39296 6 m_in[36]
port 233 nsew signal input
rlabel metal3 s 135200 40264 136000 40384 6 m_in[37]
port 234 nsew signal input
rlabel metal3 s 135200 41216 136000 41336 6 m_in[38]
port 235 nsew signal input
rlabel metal3 s 135200 42304 136000 42424 6 m_in[39]
port 236 nsew signal input
rlabel metal3 s 135200 5448 136000 5568 6 m_in[3]
port 237 nsew signal input
rlabel metal3 s 135200 43256 136000 43376 6 m_in[40]
port 238 nsew signal input
rlabel metal3 s 135200 44344 136000 44464 6 m_in[41]
port 239 nsew signal input
rlabel metal3 s 135200 45296 136000 45416 6 m_in[42]
port 240 nsew signal input
rlabel metal3 s 135200 46384 136000 46504 6 m_in[43]
port 241 nsew signal input
rlabel metal3 s 135200 47336 136000 47456 6 m_in[44]
port 242 nsew signal input
rlabel metal3 s 135200 48424 136000 48544 6 m_in[45]
port 243 nsew signal input
rlabel metal3 s 135200 49376 136000 49496 6 m_in[46]
port 244 nsew signal input
rlabel metal3 s 135200 50464 136000 50584 6 m_in[47]
port 245 nsew signal input
rlabel metal3 s 135200 51416 136000 51536 6 m_in[48]
port 246 nsew signal input
rlabel metal3 s 135200 52504 136000 52624 6 m_in[49]
port 247 nsew signal input
rlabel metal3 s 135200 6536 136000 6656 6 m_in[4]
port 248 nsew signal input
rlabel metal3 s 135200 53456 136000 53576 6 m_in[50]
port 249 nsew signal input
rlabel metal3 s 135200 54544 136000 54664 6 m_in[51]
port 250 nsew signal input
rlabel metal3 s 135200 55632 136000 55752 6 m_in[52]
port 251 nsew signal input
rlabel metal3 s 135200 56584 136000 56704 6 m_in[53]
port 252 nsew signal input
rlabel metal3 s 135200 57672 136000 57792 6 m_in[54]
port 253 nsew signal input
rlabel metal3 s 135200 58624 136000 58744 6 m_in[55]
port 254 nsew signal input
rlabel metal3 s 135200 59712 136000 59832 6 m_in[56]
port 255 nsew signal input
rlabel metal3 s 135200 60664 136000 60784 6 m_in[57]
port 256 nsew signal input
rlabel metal3 s 135200 61752 136000 61872 6 m_in[58]
port 257 nsew signal input
rlabel metal3 s 135200 62704 136000 62824 6 m_in[59]
port 258 nsew signal input
rlabel metal3 s 135200 7488 136000 7608 6 m_in[5]
port 259 nsew signal input
rlabel metal3 s 135200 63792 136000 63912 6 m_in[60]
port 260 nsew signal input
rlabel metal3 s 135200 64744 136000 64864 6 m_in[61]
port 261 nsew signal input
rlabel metal3 s 135200 65832 136000 65952 6 m_in[62]
port 262 nsew signal input
rlabel metal3 s 135200 66784 136000 66904 6 m_in[63]
port 263 nsew signal input
rlabel metal3 s 135200 67872 136000 67992 6 m_in[64]
port 264 nsew signal input
rlabel metal3 s 135200 68824 136000 68944 6 m_in[65]
port 265 nsew signal input
rlabel metal3 s 135200 69912 136000 70032 6 m_in[66]
port 266 nsew signal input
rlabel metal3 s 135200 70864 136000 70984 6 m_in[67]
port 267 nsew signal input
rlabel metal3 s 135200 71952 136000 72072 6 m_in[68]
port 268 nsew signal input
rlabel metal3 s 135200 72904 136000 73024 6 m_in[69]
port 269 nsew signal input
rlabel metal3 s 135200 8576 136000 8696 6 m_in[6]
port 270 nsew signal input
rlabel metal3 s 135200 73992 136000 74112 6 m_in[70]
port 271 nsew signal input
rlabel metal3 s 135200 74944 136000 75064 6 m_in[71]
port 272 nsew signal input
rlabel metal3 s 135200 76032 136000 76152 6 m_in[72]
port 273 nsew signal input
rlabel metal3 s 135200 76984 136000 77104 6 m_in[73]
port 274 nsew signal input
rlabel metal3 s 135200 78072 136000 78192 6 m_in[74]
port 275 nsew signal input
rlabel metal3 s 135200 79024 136000 79144 6 m_in[75]
port 276 nsew signal input
rlabel metal3 s 135200 80112 136000 80232 6 m_in[76]
port 277 nsew signal input
rlabel metal3 s 135200 81064 136000 81184 6 m_in[77]
port 278 nsew signal input
rlabel metal3 s 135200 82152 136000 82272 6 m_in[78]
port 279 nsew signal input
rlabel metal3 s 135200 83240 136000 83360 6 m_in[79]
port 280 nsew signal input
rlabel metal3 s 135200 9528 136000 9648 6 m_in[7]
port 281 nsew signal input
rlabel metal3 s 135200 84192 136000 84312 6 m_in[80]
port 282 nsew signal input
rlabel metal3 s 135200 85280 136000 85400 6 m_in[81]
port 283 nsew signal input
rlabel metal3 s 135200 86232 136000 86352 6 m_in[82]
port 284 nsew signal input
rlabel metal3 s 135200 87320 136000 87440 6 m_in[83]
port 285 nsew signal input
rlabel metal3 s 135200 88272 136000 88392 6 m_in[84]
port 286 nsew signal input
rlabel metal3 s 135200 89360 136000 89480 6 m_in[85]
port 287 nsew signal input
rlabel metal3 s 135200 90312 136000 90432 6 m_in[86]
port 288 nsew signal input
rlabel metal3 s 135200 91400 136000 91520 6 m_in[87]
port 289 nsew signal input
rlabel metal3 s 135200 92352 136000 92472 6 m_in[88]
port 290 nsew signal input
rlabel metal3 s 135200 93440 136000 93560 6 m_in[89]
port 291 nsew signal input
rlabel metal3 s 135200 10616 136000 10736 6 m_in[8]
port 292 nsew signal input
rlabel metal3 s 135200 94392 136000 94512 6 m_in[90]
port 293 nsew signal input
rlabel metal3 s 135200 95480 136000 95600 6 m_in[91]
port 294 nsew signal input
rlabel metal3 s 135200 96432 136000 96552 6 m_in[92]
port 295 nsew signal input
rlabel metal3 s 135200 97520 136000 97640 6 m_in[93]
port 296 nsew signal input
rlabel metal3 s 135200 98472 136000 98592 6 m_in[94]
port 297 nsew signal input
rlabel metal3 s 135200 99560 136000 99680 6 m_in[95]
port 298 nsew signal input
rlabel metal3 s 135200 100512 136000 100632 6 m_in[96]
port 299 nsew signal input
rlabel metal3 s 135200 101600 136000 101720 6 m_in[97]
port 300 nsew signal input
rlabel metal3 s 135200 102552 136000 102672 6 m_in[98]
port 301 nsew signal input
rlabel metal3 s 135200 103640 136000 103760 6 m_in[99]
port 302 nsew signal input
rlabel metal3 s 135200 11568 136000 11688 6 m_in[9]
port 303 nsew signal input
rlabel metal3 s 135200 1368 136000 1488 6 rst
port 304 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 stall_in
port 305 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 stall_out
port 306 nsew signal output
rlabel metal2 s 386 135200 442 136000 6 wishbone_in[0]
port 307 nsew signal input
rlabel metal2 s 8206 135200 8262 136000 6 wishbone_in[10]
port 308 nsew signal input
rlabel metal2 s 8942 135200 8998 136000 6 wishbone_in[11]
port 309 nsew signal input
rlabel metal2 s 9770 135200 9826 136000 6 wishbone_in[12]
port 310 nsew signal input
rlabel metal2 s 10598 135200 10654 136000 6 wishbone_in[13]
port 311 nsew signal input
rlabel metal2 s 11334 135200 11390 136000 6 wishbone_in[14]
port 312 nsew signal input
rlabel metal2 s 12162 135200 12218 136000 6 wishbone_in[15]
port 313 nsew signal input
rlabel metal2 s 12898 135200 12954 136000 6 wishbone_in[16]
port 314 nsew signal input
rlabel metal2 s 13726 135200 13782 136000 6 wishbone_in[17]
port 315 nsew signal input
rlabel metal2 s 14462 135200 14518 136000 6 wishbone_in[18]
port 316 nsew signal input
rlabel metal2 s 15290 135200 15346 136000 6 wishbone_in[19]
port 317 nsew signal input
rlabel metal2 s 1122 135200 1178 136000 6 wishbone_in[1]
port 318 nsew signal input
rlabel metal2 s 16026 135200 16082 136000 6 wishbone_in[20]
port 319 nsew signal input
rlabel metal2 s 16854 135200 16910 136000 6 wishbone_in[21]
port 320 nsew signal input
rlabel metal2 s 17590 135200 17646 136000 6 wishbone_in[22]
port 321 nsew signal input
rlabel metal2 s 18418 135200 18474 136000 6 wishbone_in[23]
port 322 nsew signal input
rlabel metal2 s 19246 135200 19302 136000 6 wishbone_in[24]
port 323 nsew signal input
rlabel metal2 s 19982 135200 20038 136000 6 wishbone_in[25]
port 324 nsew signal input
rlabel metal2 s 20810 135200 20866 136000 6 wishbone_in[26]
port 325 nsew signal input
rlabel metal2 s 21546 135200 21602 136000 6 wishbone_in[27]
port 326 nsew signal input
rlabel metal2 s 22374 135200 22430 136000 6 wishbone_in[28]
port 327 nsew signal input
rlabel metal2 s 23110 135200 23166 136000 6 wishbone_in[29]
port 328 nsew signal input
rlabel metal2 s 1950 135200 2006 136000 6 wishbone_in[2]
port 329 nsew signal input
rlabel metal2 s 23938 135200 23994 136000 6 wishbone_in[30]
port 330 nsew signal input
rlabel metal2 s 24674 135200 24730 136000 6 wishbone_in[31]
port 331 nsew signal input
rlabel metal2 s 25502 135200 25558 136000 6 wishbone_in[32]
port 332 nsew signal input
rlabel metal2 s 26238 135200 26294 136000 6 wishbone_in[33]
port 333 nsew signal input
rlabel metal2 s 27066 135200 27122 136000 6 wishbone_in[34]
port 334 nsew signal input
rlabel metal2 s 27894 135200 27950 136000 6 wishbone_in[35]
port 335 nsew signal input
rlabel metal2 s 28630 135200 28686 136000 6 wishbone_in[36]
port 336 nsew signal input
rlabel metal2 s 29458 135200 29514 136000 6 wishbone_in[37]
port 337 nsew signal input
rlabel metal2 s 30194 135200 30250 136000 6 wishbone_in[38]
port 338 nsew signal input
rlabel metal2 s 31022 135200 31078 136000 6 wishbone_in[39]
port 339 nsew signal input
rlabel metal2 s 2686 135200 2742 136000 6 wishbone_in[3]
port 340 nsew signal input
rlabel metal2 s 31758 135200 31814 136000 6 wishbone_in[40]
port 341 nsew signal input
rlabel metal2 s 32586 135200 32642 136000 6 wishbone_in[41]
port 342 nsew signal input
rlabel metal2 s 33322 135200 33378 136000 6 wishbone_in[42]
port 343 nsew signal input
rlabel metal2 s 34150 135200 34206 136000 6 wishbone_in[43]
port 344 nsew signal input
rlabel metal2 s 34886 135200 34942 136000 6 wishbone_in[44]
port 345 nsew signal input
rlabel metal2 s 35714 135200 35770 136000 6 wishbone_in[45]
port 346 nsew signal input
rlabel metal2 s 36450 135200 36506 136000 6 wishbone_in[46]
port 347 nsew signal input
rlabel metal2 s 37278 135200 37334 136000 6 wishbone_in[47]
port 348 nsew signal input
rlabel metal2 s 38106 135200 38162 136000 6 wishbone_in[48]
port 349 nsew signal input
rlabel metal2 s 38842 135200 38898 136000 6 wishbone_in[49]
port 350 nsew signal input
rlabel metal2 s 3514 135200 3570 136000 6 wishbone_in[4]
port 351 nsew signal input
rlabel metal2 s 39670 135200 39726 136000 6 wishbone_in[50]
port 352 nsew signal input
rlabel metal2 s 40406 135200 40462 136000 6 wishbone_in[51]
port 353 nsew signal input
rlabel metal2 s 41234 135200 41290 136000 6 wishbone_in[52]
port 354 nsew signal input
rlabel metal2 s 41970 135200 42026 136000 6 wishbone_in[53]
port 355 nsew signal input
rlabel metal2 s 42798 135200 42854 136000 6 wishbone_in[54]
port 356 nsew signal input
rlabel metal2 s 43534 135200 43590 136000 6 wishbone_in[55]
port 357 nsew signal input
rlabel metal2 s 44362 135200 44418 136000 6 wishbone_in[56]
port 358 nsew signal input
rlabel metal2 s 45098 135200 45154 136000 6 wishbone_in[57]
port 359 nsew signal input
rlabel metal2 s 45926 135200 45982 136000 6 wishbone_in[58]
port 360 nsew signal input
rlabel metal2 s 46754 135200 46810 136000 6 wishbone_in[59]
port 361 nsew signal input
rlabel metal2 s 4250 135200 4306 136000 6 wishbone_in[5]
port 362 nsew signal input
rlabel metal2 s 47490 135200 47546 136000 6 wishbone_in[60]
port 363 nsew signal input
rlabel metal2 s 48318 135200 48374 136000 6 wishbone_in[61]
port 364 nsew signal input
rlabel metal2 s 49054 135200 49110 136000 6 wishbone_in[62]
port 365 nsew signal input
rlabel metal2 s 49882 135200 49938 136000 6 wishbone_in[63]
port 366 nsew signal input
rlabel metal2 s 50618 135200 50674 136000 6 wishbone_in[64]
port 367 nsew signal input
rlabel metal2 s 51446 135200 51502 136000 6 wishbone_in[65]
port 368 nsew signal input
rlabel metal2 s 5078 135200 5134 136000 6 wishbone_in[6]
port 369 nsew signal input
rlabel metal2 s 5814 135200 5870 136000 6 wishbone_in[7]
port 370 nsew signal input
rlabel metal2 s 6642 135200 6698 136000 6 wishbone_in[8]
port 371 nsew signal input
rlabel metal2 s 7378 135200 7434 136000 6 wishbone_in[9]
port 372 nsew signal input
rlabel metal2 s 52182 135200 52238 136000 6 wishbone_out[0]
port 373 nsew signal output
rlabel metal2 s 130842 135200 130898 136000 6 wishbone_out[100]
port 374 nsew signal output
rlabel metal2 s 131578 135200 131634 136000 6 wishbone_out[101]
port 375 nsew signal output
rlabel metal2 s 132406 135200 132462 136000 6 wishbone_out[102]
port 376 nsew signal output
rlabel metal2 s 133142 135200 133198 136000 6 wishbone_out[103]
port 377 nsew signal output
rlabel metal2 s 133970 135200 134026 136000 6 wishbone_out[104]
port 378 nsew signal output
rlabel metal2 s 134706 135200 134762 136000 6 wishbone_out[105]
port 379 nsew signal output
rlabel metal2 s 135534 135200 135590 136000 6 wishbone_out[106]
port 380 nsew signal output
rlabel metal2 s 60094 135200 60150 136000 6 wishbone_out[10]
port 381 nsew signal output
rlabel metal2 s 60830 135200 60886 136000 6 wishbone_out[11]
port 382 nsew signal output
rlabel metal2 s 61658 135200 61714 136000 6 wishbone_out[12]
port 383 nsew signal output
rlabel metal2 s 62394 135200 62450 136000 6 wishbone_out[13]
port 384 nsew signal output
rlabel metal2 s 63222 135200 63278 136000 6 wishbone_out[14]
port 385 nsew signal output
rlabel metal2 s 64050 135200 64106 136000 6 wishbone_out[15]
port 386 nsew signal output
rlabel metal2 s 64786 135200 64842 136000 6 wishbone_out[16]
port 387 nsew signal output
rlabel metal2 s 65614 135200 65670 136000 6 wishbone_out[17]
port 388 nsew signal output
rlabel metal2 s 66350 135200 66406 136000 6 wishbone_out[18]
port 389 nsew signal output
rlabel metal2 s 67178 135200 67234 136000 6 wishbone_out[19]
port 390 nsew signal output
rlabel metal2 s 53010 135200 53066 136000 6 wishbone_out[1]
port 391 nsew signal output
rlabel metal2 s 67914 135200 67970 136000 6 wishbone_out[20]
port 392 nsew signal output
rlabel metal2 s 68742 135200 68798 136000 6 wishbone_out[21]
port 393 nsew signal output
rlabel metal2 s 69478 135200 69534 136000 6 wishbone_out[22]
port 394 nsew signal output
rlabel metal2 s 70306 135200 70362 136000 6 wishbone_out[23]
port 395 nsew signal output
rlabel metal2 s 71042 135200 71098 136000 6 wishbone_out[24]
port 396 nsew signal output
rlabel metal2 s 71870 135200 71926 136000 6 wishbone_out[25]
port 397 nsew signal output
rlabel metal2 s 72606 135200 72662 136000 6 wishbone_out[26]
port 398 nsew signal output
rlabel metal2 s 73434 135200 73490 136000 6 wishbone_out[27]
port 399 nsew signal output
rlabel metal2 s 74262 135200 74318 136000 6 wishbone_out[28]
port 400 nsew signal output
rlabel metal2 s 74998 135200 75054 136000 6 wishbone_out[29]
port 401 nsew signal output
rlabel metal2 s 53746 135200 53802 136000 6 wishbone_out[2]
port 402 nsew signal output
rlabel metal2 s 75826 135200 75882 136000 6 wishbone_out[30]
port 403 nsew signal output
rlabel metal2 s 76562 135200 76618 136000 6 wishbone_out[31]
port 404 nsew signal output
rlabel metal2 s 77390 135200 77446 136000 6 wishbone_out[32]
port 405 nsew signal output
rlabel metal2 s 78126 135200 78182 136000 6 wishbone_out[33]
port 406 nsew signal output
rlabel metal2 s 78954 135200 79010 136000 6 wishbone_out[34]
port 407 nsew signal output
rlabel metal2 s 79690 135200 79746 136000 6 wishbone_out[35]
port 408 nsew signal output
rlabel metal2 s 80518 135200 80574 136000 6 wishbone_out[36]
port 409 nsew signal output
rlabel metal2 s 81254 135200 81310 136000 6 wishbone_out[37]
port 410 nsew signal output
rlabel metal2 s 82082 135200 82138 136000 6 wishbone_out[38]
port 411 nsew signal output
rlabel metal2 s 82910 135200 82966 136000 6 wishbone_out[39]
port 412 nsew signal output
rlabel metal2 s 54574 135200 54630 136000 6 wishbone_out[3]
port 413 nsew signal output
rlabel metal2 s 83646 135200 83702 136000 6 wishbone_out[40]
port 414 nsew signal output
rlabel metal2 s 84474 135200 84530 136000 6 wishbone_out[41]
port 415 nsew signal output
rlabel metal2 s 85210 135200 85266 136000 6 wishbone_out[42]
port 416 nsew signal output
rlabel metal2 s 86038 135200 86094 136000 6 wishbone_out[43]
port 417 nsew signal output
rlabel metal2 s 86774 135200 86830 136000 6 wishbone_out[44]
port 418 nsew signal output
rlabel metal2 s 87602 135200 87658 136000 6 wishbone_out[45]
port 419 nsew signal output
rlabel metal2 s 88338 135200 88394 136000 6 wishbone_out[46]
port 420 nsew signal output
rlabel metal2 s 89166 135200 89222 136000 6 wishbone_out[47]
port 421 nsew signal output
rlabel metal2 s 89902 135200 89958 136000 6 wishbone_out[48]
port 422 nsew signal output
rlabel metal2 s 90730 135200 90786 136000 6 wishbone_out[49]
port 423 nsew signal output
rlabel metal2 s 55402 135200 55458 136000 6 wishbone_out[4]
port 424 nsew signal output
rlabel metal2 s 91558 135200 91614 136000 6 wishbone_out[50]
port 425 nsew signal output
rlabel metal2 s 92294 135200 92350 136000 6 wishbone_out[51]
port 426 nsew signal output
rlabel metal2 s 93122 135200 93178 136000 6 wishbone_out[52]
port 427 nsew signal output
rlabel metal2 s 93858 135200 93914 136000 6 wishbone_out[53]
port 428 nsew signal output
rlabel metal2 s 94686 135200 94742 136000 6 wishbone_out[54]
port 429 nsew signal output
rlabel metal2 s 95422 135200 95478 136000 6 wishbone_out[55]
port 430 nsew signal output
rlabel metal2 s 96250 135200 96306 136000 6 wishbone_out[56]
port 431 nsew signal output
rlabel metal2 s 96986 135200 97042 136000 6 wishbone_out[57]
port 432 nsew signal output
rlabel metal2 s 97814 135200 97870 136000 6 wishbone_out[58]
port 433 nsew signal output
rlabel metal2 s 98550 135200 98606 136000 6 wishbone_out[59]
port 434 nsew signal output
rlabel metal2 s 56138 135200 56194 136000 6 wishbone_out[5]
port 435 nsew signal output
rlabel metal2 s 99378 135200 99434 136000 6 wishbone_out[60]
port 436 nsew signal output
rlabel metal2 s 100206 135200 100262 136000 6 wishbone_out[61]
port 437 nsew signal output
rlabel metal2 s 100942 135200 100998 136000 6 wishbone_out[62]
port 438 nsew signal output
rlabel metal2 s 101770 135200 101826 136000 6 wishbone_out[63]
port 439 nsew signal output
rlabel metal2 s 102506 135200 102562 136000 6 wishbone_out[64]
port 440 nsew signal output
rlabel metal2 s 103334 135200 103390 136000 6 wishbone_out[65]
port 441 nsew signal output
rlabel metal2 s 104070 135200 104126 136000 6 wishbone_out[66]
port 442 nsew signal output
rlabel metal2 s 104898 135200 104954 136000 6 wishbone_out[67]
port 443 nsew signal output
rlabel metal2 s 105634 135200 105690 136000 6 wishbone_out[68]
port 444 nsew signal output
rlabel metal2 s 106462 135200 106518 136000 6 wishbone_out[69]
port 445 nsew signal output
rlabel metal2 s 56966 135200 57022 136000 6 wishbone_out[6]
port 446 nsew signal output
rlabel metal2 s 107198 135200 107254 136000 6 wishbone_out[70]
port 447 nsew signal output
rlabel metal2 s 108026 135200 108082 136000 6 wishbone_out[71]
port 448 nsew signal output
rlabel metal2 s 108762 135200 108818 136000 6 wishbone_out[72]
port 449 nsew signal output
rlabel metal2 s 109590 135200 109646 136000 6 wishbone_out[73]
port 450 nsew signal output
rlabel metal2 s 110418 135200 110474 136000 6 wishbone_out[74]
port 451 nsew signal output
rlabel metal2 s 111154 135200 111210 136000 6 wishbone_out[75]
port 452 nsew signal output
rlabel metal2 s 111982 135200 112038 136000 6 wishbone_out[76]
port 453 nsew signal output
rlabel metal2 s 112718 135200 112774 136000 6 wishbone_out[77]
port 454 nsew signal output
rlabel metal2 s 113546 135200 113602 136000 6 wishbone_out[78]
port 455 nsew signal output
rlabel metal2 s 114282 135200 114338 136000 6 wishbone_out[79]
port 456 nsew signal output
rlabel metal2 s 57702 135200 57758 136000 6 wishbone_out[7]
port 457 nsew signal output
rlabel metal2 s 115110 135200 115166 136000 6 wishbone_out[80]
port 458 nsew signal output
rlabel metal2 s 115846 135200 115902 136000 6 wishbone_out[81]
port 459 nsew signal output
rlabel metal2 s 116674 135200 116730 136000 6 wishbone_out[82]
port 460 nsew signal output
rlabel metal2 s 117410 135200 117466 136000 6 wishbone_out[83]
port 461 nsew signal output
rlabel metal2 s 118238 135200 118294 136000 6 wishbone_out[84]
port 462 nsew signal output
rlabel metal2 s 119066 135200 119122 136000 6 wishbone_out[85]
port 463 nsew signal output
rlabel metal2 s 119802 135200 119858 136000 6 wishbone_out[86]
port 464 nsew signal output
rlabel metal2 s 120630 135200 120686 136000 6 wishbone_out[87]
port 465 nsew signal output
rlabel metal2 s 121366 135200 121422 136000 6 wishbone_out[88]
port 466 nsew signal output
rlabel metal2 s 122194 135200 122250 136000 6 wishbone_out[89]
port 467 nsew signal output
rlabel metal2 s 58530 135200 58586 136000 6 wishbone_out[8]
port 468 nsew signal output
rlabel metal2 s 122930 135200 122986 136000 6 wishbone_out[90]
port 469 nsew signal output
rlabel metal2 s 123758 135200 123814 136000 6 wishbone_out[91]
port 470 nsew signal output
rlabel metal2 s 124494 135200 124550 136000 6 wishbone_out[92]
port 471 nsew signal output
rlabel metal2 s 125322 135200 125378 136000 6 wishbone_out[93]
port 472 nsew signal output
rlabel metal2 s 126058 135200 126114 136000 6 wishbone_out[94]
port 473 nsew signal output
rlabel metal2 s 126886 135200 126942 136000 6 wishbone_out[95]
port 474 nsew signal output
rlabel metal2 s 127714 135200 127770 136000 6 wishbone_out[96]
port 475 nsew signal output
rlabel metal2 s 128450 135200 128506 136000 6 wishbone_out[97]
port 476 nsew signal output
rlabel metal2 s 129278 135200 129334 136000 6 wishbone_out[98]
port 477 nsew signal output
rlabel metal2 s 130014 135200 130070 136000 6 wishbone_out[99]
port 478 nsew signal output
rlabel metal2 s 59266 135200 59322 136000 6 wishbone_out[9]
port 479 nsew signal output
rlabel metal4 s 127088 2128 127408 133872 6 vccd1
port 480 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 133872 6 vccd1
port 481 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 133872 6 vccd1
port 482 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 133872 6 vccd1
port 483 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 133872 6 vccd1
port 484 nsew power bidirectional
rlabel metal4 s 111728 2128 112048 133872 6 vssd1
port 485 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 133872 6 vssd1
port 486 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 133872 6 vssd1
port 487 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 133872 6 vssd1
port 488 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 136000 136000
string LEFview TRUE
string GDS_FILE /project/openlane/icache/runs/icache/results/magic/icache.gds
string GDS_END 64682064
string GDS_START 314026
<< end >>

