magic
tech sky130A
magscale 1 2
timestamp 1611902910
<< nwell >>
rect 1066 137361 209591 137371
rect 1066 136815 558846 137361
rect 1066 136805 132127 136815
rect 1066 136273 18691 136283
rect 1066 135727 558846 136273
rect 1066 135717 35067 135727
rect 1066 135185 24119 135195
rect 1066 134639 558846 135185
rect 1066 134629 11239 134639
rect 1066 134097 49787 134107
rect 1066 133551 558846 134097
rect 1066 133541 29455 133551
rect 1066 133009 33043 133019
rect 1066 132463 558846 133009
rect 1066 132453 27431 132463
rect 1066 131921 128171 131931
rect 1066 131375 558846 131921
rect 1066 131365 36079 131375
rect 1066 130833 143075 130843
rect 1066 130287 558846 130833
rect 1066 130277 40679 130287
rect 1066 129745 74903 129755
rect 1066 129199 558846 129745
rect 1066 129189 23843 129199
rect 1066 128657 107379 128667
rect 1066 128111 558846 128657
rect 1066 128101 69015 128111
rect 1066 127569 94039 127579
rect 1066 127023 558846 127569
rect 1066 127013 23843 127023
rect 1066 126481 46015 126491
rect 1066 125935 558846 126481
rect 1066 125925 38103 125935
rect 1066 125393 34883 125403
rect 1066 124847 558846 125393
rect 1066 124837 36263 124847
rect 1066 124305 16943 124315
rect 1066 123759 558846 124305
rect 1066 123749 50339 123759
rect 1066 123217 15471 123227
rect 1066 122671 558846 123217
rect 1066 122661 33135 122671
rect 1066 122129 21083 122139
rect 1066 121583 558846 122129
rect 1066 121573 46291 121583
rect 1066 121041 21083 121051
rect 1066 120495 558846 121041
rect 1066 120485 44451 120495
rect 1066 119953 40127 119963
rect 1066 119407 558846 119953
rect 1066 119397 37735 119407
rect 1066 118865 12159 118875
rect 1066 118319 558846 118865
rect 1066 118309 16851 118319
rect 1066 117777 44543 117787
rect 1066 117231 558846 117777
rect 1066 117221 57515 117231
rect 1066 116689 35711 116699
rect 1066 116143 558846 116689
rect 1066 116133 8203 116143
rect 1066 115601 21083 115611
rect 1066 115055 558846 115601
rect 1066 115045 29455 115055
rect 1066 114513 25315 114523
rect 1066 113967 558846 114513
rect 1066 113957 25223 113967
rect 1066 113425 42151 113435
rect 1066 112879 558846 113425
rect 1066 112869 33043 112879
rect 1066 112337 61287 112347
rect 1066 111791 558846 112337
rect 1066 111781 23843 111791
rect 1066 111249 18231 111259
rect 1066 110703 558846 111249
rect 1066 110693 72327 110703
rect 1066 110161 43715 110171
rect 1066 109615 558846 110161
rect 1066 109605 28075 109615
rect 1066 109073 84747 109083
rect 1066 108527 558846 109073
rect 1066 108517 24947 108527
rect 1066 107985 58803 107995
rect 1066 107439 558846 107985
rect 1066 107429 22371 107439
rect 1066 106897 100387 106907
rect 1066 106351 558846 106897
rect 1066 106341 20255 106351
rect 1066 105809 45095 105819
rect 1066 105263 558846 105809
rect 1066 105253 88335 105263
rect 1066 104721 15471 104731
rect 1066 104175 558846 104721
rect 1066 104165 37827 104175
rect 1066 103633 21635 103643
rect 1066 103087 558846 103633
rect 1066 103077 29455 103087
rect 1066 102545 40863 102555
rect 1066 101999 558846 102545
rect 1066 101989 29915 101999
rect 1066 101457 22647 101467
rect 1066 100911 558846 101457
rect 1066 100901 63403 100911
rect 1066 100369 82815 100379
rect 1066 99823 558846 100369
rect 1066 99813 44911 99823
rect 1066 99281 49143 99291
rect 1066 98735 558846 99281
rect 1066 98725 74351 98735
rect 1066 98193 22923 98203
rect 1066 97647 558846 98193
rect 1066 97637 18599 97647
rect 1066 97105 16943 97115
rect 1066 96559 558846 97105
rect 1066 96549 96799 96559
rect 1066 96017 46015 96027
rect 1066 95471 558846 96017
rect 1066 95461 27247 95471
rect 1066 94929 34699 94939
rect 1066 94383 558846 94929
rect 1066 94373 16299 94383
rect 1066 93841 32307 93851
rect 1066 93295 558846 93841
rect 1066 93285 35895 93295
rect 1066 92753 21543 92763
rect 1066 92207 558846 92753
rect 1066 92197 102411 92207
rect 1066 91665 94039 91675
rect 1066 91119 558846 91665
rect 1066 91109 18231 91119
rect 1066 90577 24395 90587
rect 1066 90031 558846 90577
rect 1066 90021 19427 90031
rect 1066 89489 24395 89499
rect 1066 88943 558846 89489
rect 1066 88933 52547 88943
rect 1066 88401 11423 88411
rect 1066 87855 558846 88401
rect 1066 87845 20531 87855
rect 1066 87313 18599 87323
rect 1066 86767 558846 87313
rect 1066 86757 72051 86767
rect 1066 86225 25315 86235
rect 1066 85679 558846 86225
rect 1066 85669 18231 85679
rect 1066 85137 25315 85147
rect 1066 84591 558846 85137
rect 1066 84581 14091 84591
rect 1066 84049 19059 84059
rect 1066 83503 558846 84049
rect 1066 83493 21083 83503
rect 1066 82961 24303 82971
rect 1066 82415 558846 82961
rect 1066 82405 59999 82415
rect 1066 81873 12895 81883
rect 1066 81327 558846 81873
rect 1066 81317 15379 81327
rect 1066 80785 18967 80795
rect 1066 80239 558846 80785
rect 1066 80229 26327 80239
rect 1066 79697 43531 79707
rect 1066 79151 558846 79697
rect 1066 79141 63311 79151
rect 1066 78609 98271 78619
rect 1066 78063 558846 78609
rect 1066 78053 98363 78063
rect 1066 77521 199103 77531
rect 1066 76975 558846 77521
rect 1066 76965 165707 76975
rect 1066 76433 15471 76443
rect 1066 75887 558846 76433
rect 1066 75877 33319 75887
rect 1066 75345 18691 75355
rect 1066 74799 558846 75345
rect 1066 74789 19703 74799
rect 1066 74257 12435 74267
rect 1066 73711 558846 74257
rect 1066 73701 7099 73711
rect 1066 73169 119339 73179
rect 1066 72623 558846 73169
rect 1066 72613 29639 72623
rect 1066 72081 21083 72091
rect 1066 71535 558846 72081
rect 1066 71525 20715 71535
rect 1066 70993 28627 71003
rect 1066 70447 558846 70993
rect 1066 70437 12619 70447
rect 1066 69905 16943 69915
rect 1066 69359 558846 69905
rect 1066 69349 22279 69359
rect 1066 68817 21083 68827
rect 1066 68271 558846 68817
rect 1066 68261 80699 68271
rect 1066 67729 16391 67739
rect 1066 67183 558846 67729
rect 1066 67173 29915 67183
rect 1066 66641 23107 66651
rect 1066 66095 558846 66641
rect 1066 66085 11239 66095
rect 1066 65553 28903 65563
rect 1066 65007 558846 65553
rect 1066 64997 29455 65007
rect 1066 64465 7007 64475
rect 1066 63919 558846 64465
rect 1066 63909 23843 63919
rect 1066 63377 28995 63387
rect 1066 62831 558846 63377
rect 1066 62821 21727 62831
rect 1066 62289 24211 62299
rect 1066 61743 558846 62289
rect 1066 61733 2407 61743
rect 1066 61201 229739 61211
rect 1066 60655 558846 61201
rect 1066 60645 117775 60655
rect 1066 60113 97903 60123
rect 1066 59567 558846 60113
rect 1066 59557 12803 59567
rect 1066 59025 36355 59035
rect 1066 58479 558846 59025
rect 1066 58469 3327 58479
rect 1066 57937 45923 57947
rect 1066 57391 558846 57937
rect 1066 57381 81987 57391
rect 1066 56849 24119 56859
rect 1066 56303 558846 56849
rect 1066 56293 15839 56303
rect 1066 55761 21083 55771
rect 1066 55215 558846 55761
rect 1066 55205 12803 55215
rect 1066 54673 22739 54683
rect 1066 54127 558846 54673
rect 1066 54117 59631 54127
rect 1066 53585 26695 53595
rect 1066 53039 558846 53585
rect 1066 53029 39299 53039
rect 1066 52497 23015 52507
rect 1066 51951 558846 52497
rect 1066 51941 40679 51951
rect 1066 51409 27155 51419
rect 1066 50863 558846 51409
rect 1066 50853 24579 50863
rect 1066 50321 13723 50331
rect 1066 49775 558846 50321
rect 1066 49765 14827 49775
rect 1066 49233 12527 49243
rect 1066 48687 558846 49233
rect 1066 48677 23843 48687
rect 1066 48145 9951 48155
rect 1066 47599 558846 48145
rect 1066 47589 10227 47599
rect 1066 47057 183831 47067
rect 1066 46511 558846 47057
rect 1066 46501 43163 46511
rect 1066 45969 69199 45979
rect 1066 45423 558846 45969
rect 1066 45413 33043 45423
rect 1066 44881 22555 44891
rect 1066 44335 558846 44881
rect 1066 44325 19795 44335
rect 1066 43793 18875 43803
rect 1066 43247 558846 43793
rect 1066 43237 23843 43247
rect 1066 42705 112531 42715
rect 1066 42159 558846 42705
rect 1066 42149 70671 42159
rect 1066 41617 17035 41627
rect 1066 41071 558846 41617
rect 1066 41061 18875 41071
rect 1066 40529 43807 40539
rect 1066 39983 558846 40529
rect 1066 39973 10411 39983
rect 1066 39441 25223 39451
rect 1066 38895 558846 39441
rect 1066 38885 19519 38895
rect 1066 38353 19151 38363
rect 1066 37807 558846 38353
rect 1066 37797 71867 37807
rect 1066 37265 43531 37275
rect 1066 36719 558846 37265
rect 1066 36709 78307 36719
rect 1066 36177 78307 36187
rect 1066 35631 558846 36177
rect 1066 35621 27339 35631
rect 1066 35089 8479 35099
rect 1066 34543 558846 35089
rect 1066 34533 85575 34543
rect 1066 34001 49143 34011
rect 1066 33455 558846 34001
rect 1066 33445 31571 33455
rect 1066 32913 46751 32923
rect 1066 32367 558846 32913
rect 1066 32357 8203 32367
rect 1066 31825 43531 31835
rect 1066 31279 558846 31825
rect 1066 31269 12619 31279
rect 1066 30737 38931 30747
rect 1066 30191 558846 30737
rect 1066 30181 21727 30191
rect 1066 29649 28167 29659
rect 1066 29103 558846 29649
rect 1066 29093 7007 29103
rect 1066 28561 74719 28571
rect 1066 28015 558846 28561
rect 1066 28005 22003 28015
rect 1066 27473 24855 27483
rect 1066 26927 558846 27473
rect 1066 26917 23843 26927
rect 1066 26385 13355 26395
rect 1066 25839 558846 26385
rect 1066 25829 35067 25839
rect 1066 25297 38655 25307
rect 1066 24751 558846 25297
rect 1066 24741 40679 24751
rect 1066 24209 9859 24219
rect 1066 23663 558846 24209
rect 1066 23653 18231 23663
rect 1066 23121 17311 23131
rect 1066 22575 558846 23121
rect 1066 22565 42151 22575
rect 1066 22033 21083 22043
rect 1066 21487 558846 22033
rect 1066 21477 8847 21487
rect 1066 20945 32307 20955
rect 1066 20399 558846 20945
rect 1066 20389 27523 20399
rect 1066 19857 39943 19867
rect 1066 19311 558846 19857
rect 1066 19301 29455 19311
rect 1066 18769 84931 18779
rect 1066 18223 558846 18769
rect 1066 18213 63127 18223
rect 1066 17681 11515 17691
rect 1066 17135 558846 17681
rect 1066 17125 18231 17135
rect 1066 16593 6363 16603
rect 1066 16047 558846 16593
rect 1066 16037 61747 16047
rect 1066 15505 27247 15515
rect 1066 14959 558846 15505
rect 1066 14949 9675 14959
rect 1066 14417 22739 14427
rect 1066 13871 558846 14417
rect 1066 13861 23843 13871
rect 1066 13329 7743 13339
rect 1066 12783 558846 13329
rect 1066 12773 40679 12783
rect 1066 12241 28167 12251
rect 1066 11695 558846 12241
rect 1066 11685 8663 11695
rect 1066 11153 62299 11163
rect 1066 10607 558846 11153
rect 1066 10597 2591 10607
rect 1066 10065 37919 10075
rect 1066 9519 558846 10065
rect 1066 9509 9859 9519
rect 1066 8977 18415 8987
rect 1066 8431 558846 8977
rect 1066 8421 25775 8431
rect 1066 7889 23107 7899
rect 1066 7343 558846 7889
rect 1066 7333 20071 7343
rect 1066 6801 45003 6811
rect 1066 6255 558846 6801
rect 1066 6245 48315 6255
rect 1066 5713 68095 5723
rect 1066 5167 558846 5713
rect 1066 5157 55491 5167
rect 1066 4625 114371 4635
rect 1066 4079 558846 4625
rect 1066 4069 164143 4079
rect 1066 3537 347867 3547
rect 1066 2991 558846 3537
rect 1066 2981 190179 2991
rect 1066 2138 558846 2459
<< obsli1 >>
rect 1104 1309 558808 138091
<< obsm1 >>
rect 1104 1164 558808 138100
<< metal2 >>
rect 1858 0 1914 800
rect 5630 0 5686 800
rect 9402 0 9458 800
rect 13266 0 13322 800
rect 17038 0 17094 800
rect 20902 0 20958 800
rect 24674 0 24730 800
rect 28446 0 28502 800
rect 32310 0 32366 800
rect 36082 0 36138 800
rect 39946 0 40002 800
rect 43718 0 43774 800
rect 47490 0 47546 800
rect 51354 0 51410 800
rect 55126 0 55182 800
rect 58990 0 59046 800
rect 62762 0 62818 800
rect 66534 0 66590 800
rect 70398 0 70454 800
rect 74170 0 74226 800
rect 78034 0 78090 800
rect 81806 0 81862 800
rect 85578 0 85634 800
rect 89442 0 89498 800
rect 93214 0 93270 800
rect 97078 0 97134 800
rect 100850 0 100906 800
rect 104714 0 104770 800
rect 108486 0 108542 800
rect 112258 0 112314 800
rect 116122 0 116178 800
rect 119894 0 119950 800
rect 123758 0 123814 800
rect 127530 0 127586 800
rect 131302 0 131358 800
rect 135166 0 135222 800
rect 138938 0 138994 800
rect 142802 0 142858 800
rect 146574 0 146630 800
rect 150346 0 150402 800
rect 154210 0 154266 800
rect 157982 0 158038 800
rect 161846 0 161902 800
rect 165618 0 165674 800
rect 169390 0 169446 800
rect 173254 0 173310 800
rect 177026 0 177082 800
rect 180890 0 180946 800
rect 184662 0 184718 800
rect 188526 0 188582 800
rect 192298 0 192354 800
rect 196070 0 196126 800
rect 199934 0 199990 800
rect 203706 0 203762 800
rect 207570 0 207626 800
rect 211342 0 211398 800
rect 215114 0 215170 800
rect 218978 0 219034 800
rect 222750 0 222806 800
rect 226614 0 226670 800
rect 230386 0 230442 800
rect 234158 0 234214 800
rect 238022 0 238078 800
rect 241794 0 241850 800
rect 245658 0 245714 800
rect 249430 0 249486 800
rect 253202 0 253258 800
rect 257066 0 257122 800
rect 260838 0 260894 800
rect 264702 0 264758 800
rect 268474 0 268530 800
rect 272246 0 272302 800
rect 276110 0 276166 800
rect 279882 0 279938 800
rect 283746 0 283802 800
rect 287518 0 287574 800
rect 291382 0 291438 800
rect 295154 0 295210 800
rect 298926 0 298982 800
rect 302790 0 302846 800
rect 306562 0 306618 800
rect 310426 0 310482 800
rect 314198 0 314254 800
rect 317970 0 318026 800
rect 321834 0 321890 800
rect 325606 0 325662 800
rect 329470 0 329526 800
rect 333242 0 333298 800
rect 337014 0 337070 800
rect 340878 0 340934 800
rect 344650 0 344706 800
rect 348514 0 348570 800
rect 352286 0 352342 800
rect 356058 0 356114 800
rect 359922 0 359978 800
rect 363694 0 363750 800
rect 367558 0 367614 800
rect 371330 0 371386 800
rect 375194 0 375250 800
rect 378966 0 379022 800
rect 382738 0 382794 800
rect 386602 0 386658 800
rect 390374 0 390430 800
rect 394238 0 394294 800
rect 398010 0 398066 800
rect 401782 0 401838 800
rect 405646 0 405702 800
rect 409418 0 409474 800
rect 413282 0 413338 800
rect 417054 0 417110 800
rect 420826 0 420882 800
rect 424690 0 424746 800
rect 428462 0 428518 800
rect 432326 0 432382 800
rect 436098 0 436154 800
rect 439870 0 439926 800
rect 443734 0 443790 800
rect 447506 0 447562 800
rect 451370 0 451426 800
rect 455142 0 455198 800
rect 458914 0 458970 800
rect 462778 0 462834 800
rect 466550 0 466606 800
rect 470414 0 470470 800
rect 474186 0 474242 800
rect 478050 0 478106 800
rect 481822 0 481878 800
rect 485594 0 485650 800
rect 489458 0 489514 800
rect 493230 0 493286 800
rect 497094 0 497150 800
rect 500866 0 500922 800
rect 504638 0 504694 800
rect 508502 0 508558 800
rect 512274 0 512330 800
rect 516138 0 516194 800
rect 519910 0 519966 800
rect 523682 0 523738 800
rect 527546 0 527602 800
rect 531318 0 531374 800
rect 535182 0 535238 800
rect 538954 0 539010 800
rect 542726 0 542782 800
rect 546590 0 546646 800
rect 550362 0 550418 800
rect 554226 0 554282 800
rect 557998 0 558054 800
<< obsm2 >>
rect 1860 856 558236 138106
rect 1970 800 5574 856
rect 5742 800 9346 856
rect 9514 800 13210 856
rect 13378 800 16982 856
rect 17150 800 20846 856
rect 21014 800 24618 856
rect 24786 800 28390 856
rect 28558 800 32254 856
rect 32422 800 36026 856
rect 36194 800 39890 856
rect 40058 800 43662 856
rect 43830 800 47434 856
rect 47602 800 51298 856
rect 51466 800 55070 856
rect 55238 800 58934 856
rect 59102 800 62706 856
rect 62874 800 66478 856
rect 66646 800 70342 856
rect 70510 800 74114 856
rect 74282 800 77978 856
rect 78146 800 81750 856
rect 81918 800 85522 856
rect 85690 800 89386 856
rect 89554 800 93158 856
rect 93326 800 97022 856
rect 97190 800 100794 856
rect 100962 800 104658 856
rect 104826 800 108430 856
rect 108598 800 112202 856
rect 112370 800 116066 856
rect 116234 800 119838 856
rect 120006 800 123702 856
rect 123870 800 127474 856
rect 127642 800 131246 856
rect 131414 800 135110 856
rect 135278 800 138882 856
rect 139050 800 142746 856
rect 142914 800 146518 856
rect 146686 800 150290 856
rect 150458 800 154154 856
rect 154322 800 157926 856
rect 158094 800 161790 856
rect 161958 800 165562 856
rect 165730 800 169334 856
rect 169502 800 173198 856
rect 173366 800 176970 856
rect 177138 800 180834 856
rect 181002 800 184606 856
rect 184774 800 188470 856
rect 188638 800 192242 856
rect 192410 800 196014 856
rect 196182 800 199878 856
rect 200046 800 203650 856
rect 203818 800 207514 856
rect 207682 800 211286 856
rect 211454 800 215058 856
rect 215226 800 218922 856
rect 219090 800 222694 856
rect 222862 800 226558 856
rect 226726 800 230330 856
rect 230498 800 234102 856
rect 234270 800 237966 856
rect 238134 800 241738 856
rect 241906 800 245602 856
rect 245770 800 249374 856
rect 249542 800 253146 856
rect 253314 800 257010 856
rect 257178 800 260782 856
rect 260950 800 264646 856
rect 264814 800 268418 856
rect 268586 800 272190 856
rect 272358 800 276054 856
rect 276222 800 279826 856
rect 279994 800 283690 856
rect 283858 800 287462 856
rect 287630 800 291326 856
rect 291494 800 295098 856
rect 295266 800 298870 856
rect 299038 800 302734 856
rect 302902 800 306506 856
rect 306674 800 310370 856
rect 310538 800 314142 856
rect 314310 800 317914 856
rect 318082 800 321778 856
rect 321946 800 325550 856
rect 325718 800 329414 856
rect 329582 800 333186 856
rect 333354 800 336958 856
rect 337126 800 340822 856
rect 340990 800 344594 856
rect 344762 800 348458 856
rect 348626 800 352230 856
rect 352398 800 356002 856
rect 356170 800 359866 856
rect 360034 800 363638 856
rect 363806 800 367502 856
rect 367670 800 371274 856
rect 371442 800 375138 856
rect 375306 800 378910 856
rect 379078 800 382682 856
rect 382850 800 386546 856
rect 386714 800 390318 856
rect 390486 800 394182 856
rect 394350 800 397954 856
rect 398122 800 401726 856
rect 401894 800 405590 856
rect 405758 800 409362 856
rect 409530 800 413226 856
rect 413394 800 416998 856
rect 417166 800 420770 856
rect 420938 800 424634 856
rect 424802 800 428406 856
rect 428574 800 432270 856
rect 432438 800 436042 856
rect 436210 800 439814 856
rect 439982 800 443678 856
rect 443846 800 447450 856
rect 447618 800 451314 856
rect 451482 800 455086 856
rect 455254 800 458858 856
rect 459026 800 462722 856
rect 462890 800 466494 856
rect 466662 800 470358 856
rect 470526 800 474130 856
rect 474298 800 477994 856
rect 478162 800 481766 856
rect 481934 800 485538 856
rect 485706 800 489402 856
rect 489570 800 493174 856
rect 493342 800 497038 856
rect 497206 800 500810 856
rect 500978 800 504582 856
rect 504750 800 508446 856
rect 508614 800 512218 856
rect 512386 800 516082 856
rect 516250 800 519854 856
rect 520022 800 523626 856
rect 523794 800 527490 856
rect 527658 800 531262 856
rect 531430 800 535126 856
rect 535294 800 538898 856
rect 539066 800 542670 856
rect 542838 800 546534 856
rect 546702 800 550306 856
rect 550474 800 554170 856
rect 554338 800 557942 856
rect 558110 800 558236 856
<< obsm3 >>
rect 2589 1803 558059 137733
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
rect 142448 2128 142768 137680
rect 157808 2128 158128 137680
rect 173168 2128 173488 137680
rect 188528 2128 188848 137680
rect 203888 2128 204208 137680
rect 219248 2128 219568 137680
rect 234608 2128 234928 137680
rect 249968 2128 250288 137680
rect 265328 2128 265648 137680
rect 280688 2128 281008 137680
rect 296048 2128 296368 137680
rect 311408 2128 311728 137680
rect 326768 2128 327088 137680
rect 342128 2128 342448 137680
rect 357488 2128 357808 137680
rect 372848 2128 373168 137680
rect 388208 2128 388528 137680
rect 403568 2128 403888 137680
rect 418928 2128 419248 137680
rect 434288 2128 434608 137680
rect 449648 2128 449968 137680
rect 465008 2128 465328 137680
rect 480368 2128 480688 137680
rect 495728 2128 496048 137680
rect 511088 2128 511408 137680
rect 526448 2128 526768 137680
rect 541808 2128 542128 137680
rect 557168 2128 557488 137680
<< obsm4 >>
rect 19379 2048 19488 134605
rect 19968 2048 34848 134605
rect 35328 2048 50208 134605
rect 50688 2048 65568 134605
rect 66048 2048 80928 134605
rect 81408 2048 96288 134605
rect 96768 2048 111648 134605
rect 112128 2048 127008 134605
rect 127488 2048 142368 134605
rect 142848 2048 157728 134605
rect 158208 2048 173088 134605
rect 173568 2048 188448 134605
rect 188928 2048 203808 134605
rect 204288 2048 219168 134605
rect 219648 2048 234528 134605
rect 235008 2048 249888 134605
rect 250368 2048 265248 134605
rect 265728 2048 280608 134605
rect 281088 2048 295968 134605
rect 296448 2048 311328 134605
rect 311808 2048 326688 134605
rect 327168 2048 342048 134605
rect 342528 2048 357408 134605
rect 357888 2048 372768 134605
rect 373248 2048 388128 134605
rect 388608 2048 403488 134605
rect 403968 2048 418848 134605
rect 419328 2048 434208 134605
rect 434688 2048 449568 134605
rect 450048 2048 464928 134605
rect 465408 2048 480288 134605
rect 480768 2048 495648 134605
rect 496128 2048 511008 134605
rect 511488 2048 526368 134605
rect 526848 2048 541728 134605
rect 542208 2048 543845 134605
rect 19379 1803 543845 2048
<< labels >>
rlabel metal2 s 489458 0 489514 800 6 A[0]
port 1 nsew signal input
rlabel metal2 s 493230 0 493286 800 6 A[1]
port 2 nsew signal input
rlabel metal2 s 497094 0 497150 800 6 A[2]
port 3 nsew signal input
rlabel metal2 s 500866 0 500922 800 6 A[3]
port 4 nsew signal input
rlabel metal2 s 504638 0 504694 800 6 A[4]
port 5 nsew signal input
rlabel metal2 s 508502 0 508558 800 6 A[5]
port 6 nsew signal input
rlabel metal2 s 512274 0 512330 800 6 A[6]
port 7 nsew signal input
rlabel metal2 s 516138 0 516194 800 6 A[7]
port 8 nsew signal input
rlabel metal2 s 519910 0 519966 800 6 A[8]
port 9 nsew signal input
rlabel metal2 s 523682 0 523738 800 6 CLK
port 10 nsew signal input
rlabel metal2 s 245658 0 245714 800 6 Di[0]
port 11 nsew signal input
rlabel metal2 s 283746 0 283802 800 6 Di[10]
port 12 nsew signal input
rlabel metal2 s 287518 0 287574 800 6 Di[11]
port 13 nsew signal input
rlabel metal2 s 291382 0 291438 800 6 Di[12]
port 14 nsew signal input
rlabel metal2 s 295154 0 295210 800 6 Di[13]
port 15 nsew signal input
rlabel metal2 s 298926 0 298982 800 6 Di[14]
port 16 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 Di[15]
port 17 nsew signal input
rlabel metal2 s 306562 0 306618 800 6 Di[16]
port 18 nsew signal input
rlabel metal2 s 310426 0 310482 800 6 Di[17]
port 19 nsew signal input
rlabel metal2 s 314198 0 314254 800 6 Di[18]
port 20 nsew signal input
rlabel metal2 s 317970 0 318026 800 6 Di[19]
port 21 nsew signal input
rlabel metal2 s 249430 0 249486 800 6 Di[1]
port 22 nsew signal input
rlabel metal2 s 321834 0 321890 800 6 Di[20]
port 23 nsew signal input
rlabel metal2 s 325606 0 325662 800 6 Di[21]
port 24 nsew signal input
rlabel metal2 s 329470 0 329526 800 6 Di[22]
port 25 nsew signal input
rlabel metal2 s 333242 0 333298 800 6 Di[23]
port 26 nsew signal input
rlabel metal2 s 337014 0 337070 800 6 Di[24]
port 27 nsew signal input
rlabel metal2 s 340878 0 340934 800 6 Di[25]
port 28 nsew signal input
rlabel metal2 s 344650 0 344706 800 6 Di[26]
port 29 nsew signal input
rlabel metal2 s 348514 0 348570 800 6 Di[27]
port 30 nsew signal input
rlabel metal2 s 352286 0 352342 800 6 Di[28]
port 31 nsew signal input
rlabel metal2 s 356058 0 356114 800 6 Di[29]
port 32 nsew signal input
rlabel metal2 s 253202 0 253258 800 6 Di[2]
port 33 nsew signal input
rlabel metal2 s 359922 0 359978 800 6 Di[30]
port 34 nsew signal input
rlabel metal2 s 363694 0 363750 800 6 Di[31]
port 35 nsew signal input
rlabel metal2 s 367558 0 367614 800 6 Di[32]
port 36 nsew signal input
rlabel metal2 s 371330 0 371386 800 6 Di[33]
port 37 nsew signal input
rlabel metal2 s 375194 0 375250 800 6 Di[34]
port 38 nsew signal input
rlabel metal2 s 378966 0 379022 800 6 Di[35]
port 39 nsew signal input
rlabel metal2 s 382738 0 382794 800 6 Di[36]
port 40 nsew signal input
rlabel metal2 s 386602 0 386658 800 6 Di[37]
port 41 nsew signal input
rlabel metal2 s 390374 0 390430 800 6 Di[38]
port 42 nsew signal input
rlabel metal2 s 394238 0 394294 800 6 Di[39]
port 43 nsew signal input
rlabel metal2 s 257066 0 257122 800 6 Di[3]
port 44 nsew signal input
rlabel metal2 s 398010 0 398066 800 6 Di[40]
port 45 nsew signal input
rlabel metal2 s 401782 0 401838 800 6 Di[41]
port 46 nsew signal input
rlabel metal2 s 405646 0 405702 800 6 Di[42]
port 47 nsew signal input
rlabel metal2 s 409418 0 409474 800 6 Di[43]
port 48 nsew signal input
rlabel metal2 s 413282 0 413338 800 6 Di[44]
port 49 nsew signal input
rlabel metal2 s 417054 0 417110 800 6 Di[45]
port 50 nsew signal input
rlabel metal2 s 420826 0 420882 800 6 Di[46]
port 51 nsew signal input
rlabel metal2 s 424690 0 424746 800 6 Di[47]
port 52 nsew signal input
rlabel metal2 s 428462 0 428518 800 6 Di[48]
port 53 nsew signal input
rlabel metal2 s 432326 0 432382 800 6 Di[49]
port 54 nsew signal input
rlabel metal2 s 260838 0 260894 800 6 Di[4]
port 55 nsew signal input
rlabel metal2 s 436098 0 436154 800 6 Di[50]
port 56 nsew signal input
rlabel metal2 s 439870 0 439926 800 6 Di[51]
port 57 nsew signal input
rlabel metal2 s 443734 0 443790 800 6 Di[52]
port 58 nsew signal input
rlabel metal2 s 447506 0 447562 800 6 Di[53]
port 59 nsew signal input
rlabel metal2 s 451370 0 451426 800 6 Di[54]
port 60 nsew signal input
rlabel metal2 s 455142 0 455198 800 6 Di[55]
port 61 nsew signal input
rlabel metal2 s 458914 0 458970 800 6 Di[56]
port 62 nsew signal input
rlabel metal2 s 462778 0 462834 800 6 Di[57]
port 63 nsew signal input
rlabel metal2 s 466550 0 466606 800 6 Di[58]
port 64 nsew signal input
rlabel metal2 s 470414 0 470470 800 6 Di[59]
port 65 nsew signal input
rlabel metal2 s 264702 0 264758 800 6 Di[5]
port 66 nsew signal input
rlabel metal2 s 474186 0 474242 800 6 Di[60]
port 67 nsew signal input
rlabel metal2 s 478050 0 478106 800 6 Di[61]
port 68 nsew signal input
rlabel metal2 s 481822 0 481878 800 6 Di[62]
port 69 nsew signal input
rlabel metal2 s 485594 0 485650 800 6 Di[63]
port 70 nsew signal input
rlabel metal2 s 268474 0 268530 800 6 Di[6]
port 71 nsew signal input
rlabel metal2 s 272246 0 272302 800 6 Di[7]
port 72 nsew signal input
rlabel metal2 s 276110 0 276166 800 6 Di[8]
port 73 nsew signal input
rlabel metal2 s 279882 0 279938 800 6 Di[9]
port 74 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 Do[0]
port 75 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 Do[10]
port 76 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 Do[11]
port 77 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 Do[12]
port 78 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 Do[13]
port 79 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 Do[14]
port 80 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 Do[15]
port 81 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 Do[16]
port 82 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 Do[17]
port 83 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 Do[18]
port 84 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 Do[19]
port 85 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 Do[1]
port 86 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 Do[20]
port 87 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 Do[21]
port 88 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 Do[22]
port 89 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 Do[23]
port 90 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 Do[24]
port 91 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 Do[25]
port 92 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 Do[26]
port 93 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 Do[27]
port 94 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 Do[28]
port 95 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 Do[29]
port 96 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 Do[2]
port 97 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 Do[30]
port 98 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 Do[31]
port 99 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 Do[32]
port 100 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 Do[33]
port 101 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 Do[34]
port 102 nsew signal output
rlabel metal2 s 135166 0 135222 800 6 Do[35]
port 103 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 Do[36]
port 104 nsew signal output
rlabel metal2 s 142802 0 142858 800 6 Do[37]
port 105 nsew signal output
rlabel metal2 s 146574 0 146630 800 6 Do[38]
port 106 nsew signal output
rlabel metal2 s 150346 0 150402 800 6 Do[39]
port 107 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 Do[3]
port 108 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 Do[40]
port 109 nsew signal output
rlabel metal2 s 157982 0 158038 800 6 Do[41]
port 110 nsew signal output
rlabel metal2 s 161846 0 161902 800 6 Do[42]
port 111 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 Do[43]
port 112 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 Do[44]
port 113 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 Do[45]
port 114 nsew signal output
rlabel metal2 s 177026 0 177082 800 6 Do[46]
port 115 nsew signal output
rlabel metal2 s 180890 0 180946 800 6 Do[47]
port 116 nsew signal output
rlabel metal2 s 184662 0 184718 800 6 Do[48]
port 117 nsew signal output
rlabel metal2 s 188526 0 188582 800 6 Do[49]
port 118 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 Do[4]
port 119 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 Do[50]
port 120 nsew signal output
rlabel metal2 s 196070 0 196126 800 6 Do[51]
port 121 nsew signal output
rlabel metal2 s 199934 0 199990 800 6 Do[52]
port 122 nsew signal output
rlabel metal2 s 203706 0 203762 800 6 Do[53]
port 123 nsew signal output
rlabel metal2 s 207570 0 207626 800 6 Do[54]
port 124 nsew signal output
rlabel metal2 s 211342 0 211398 800 6 Do[55]
port 125 nsew signal output
rlabel metal2 s 215114 0 215170 800 6 Do[56]
port 126 nsew signal output
rlabel metal2 s 218978 0 219034 800 6 Do[57]
port 127 nsew signal output
rlabel metal2 s 222750 0 222806 800 6 Do[58]
port 128 nsew signal output
rlabel metal2 s 226614 0 226670 800 6 Do[59]
port 129 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 Do[5]
port 130 nsew signal output
rlabel metal2 s 230386 0 230442 800 6 Do[60]
port 131 nsew signal output
rlabel metal2 s 234158 0 234214 800 6 Do[61]
port 132 nsew signal output
rlabel metal2 s 238022 0 238078 800 6 Do[62]
port 133 nsew signal output
rlabel metal2 s 241794 0 241850 800 6 Do[63]
port 134 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 Do[6]
port 135 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 Do[7]
port 136 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 Do[8]
port 137 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 Do[9]
port 138 nsew signal output
rlabel metal2 s 557998 0 558054 800 6 EN
port 139 nsew signal input
rlabel metal2 s 527546 0 527602 800 6 WE[0]
port 140 nsew signal input
rlabel metal2 s 531318 0 531374 800 6 WE[1]
port 141 nsew signal input
rlabel metal2 s 535182 0 535238 800 6 WE[2]
port 142 nsew signal input
rlabel metal2 s 538954 0 539010 800 6 WE[3]
port 143 nsew signal input
rlabel metal2 s 542726 0 542782 800 6 WE[4]
port 144 nsew signal input
rlabel metal2 s 546590 0 546646 800 6 WE[5]
port 145 nsew signal input
rlabel metal2 s 550362 0 550418 800 6 WE[6]
port 146 nsew signal input
rlabel metal2 s 554226 0 554282 800 6 WE[7]
port 147 nsew signal input
rlabel metal4 s 557168 2128 557488 137680 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 137680 6 vccd1
port 149 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 137680 6 vccd1
port 150 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 137680 6 vccd1
port 151 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 137680 6 vccd1
port 152 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 137680 6 vccd1
port 153 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 137680 6 vccd1
port 154 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 137680 6 vccd1
port 155 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 137680 6 vccd1
port 156 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 137680 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 137680 6 vccd1
port 158 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 137680 6 vccd1
port 159 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 137680 6 vccd1
port 160 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 137680 6 vccd1
port 161 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 162 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 163 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 164 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 165 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 166 nsew power bidirectional
rlabel metal4 s 541808 2128 542128 137680 6 vssd1
port 167 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 137680 6 vssd1
port 168 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 137680 6 vssd1
port 169 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 137680 6 vssd1
port 170 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 137680 6 vssd1
port 171 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 137680 6 vssd1
port 172 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 137680 6 vssd1
port 173 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 137680 6 vssd1
port 174 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 137680 6 vssd1
port 175 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 137680 6 vssd1
port 176 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 137680 6 vssd1
port 177 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 137680 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 137680 6 vssd1
port 179 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 137680 6 vssd1
port 180 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 181 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 182 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 183 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 184 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 560000 140000
string LEFview TRUE
string GDS_FILE /project/openlane/RAM_512x64/runs/RAM_512x64/results/magic/RAM_512x64.gds
string GDS_END 298454472
string GDS_START 192796
<< end >>

