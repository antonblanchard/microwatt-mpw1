magic
tech sky130A
magscale 1 2
timestamp 1612123974
<< obsli1 >>
rect 1104 2159 219023 217617
<< obsm1 >>
rect 1104 2128 219406 218408
<< metal2 >>
rect 478 219200 534 220000
rect 1490 219200 1546 220000
rect 2502 219200 2558 220000
rect 3514 219200 3570 220000
rect 4526 219200 4582 220000
rect 5538 219200 5594 220000
rect 6550 219200 6606 220000
rect 7562 219200 7618 220000
rect 8574 219200 8630 220000
rect 9586 219200 9642 220000
rect 10598 219200 10654 220000
rect 11610 219200 11666 220000
rect 12622 219200 12678 220000
rect 13634 219200 13690 220000
rect 14646 219200 14702 220000
rect 15658 219200 15714 220000
rect 16670 219200 16726 220000
rect 17682 219200 17738 220000
rect 18694 219200 18750 220000
rect 19706 219200 19762 220000
rect 20718 219200 20774 220000
rect 21730 219200 21786 220000
rect 22742 219200 22798 220000
rect 23754 219200 23810 220000
rect 24766 219200 24822 220000
rect 25778 219200 25834 220000
rect 26790 219200 26846 220000
rect 27802 219200 27858 220000
rect 28814 219200 28870 220000
rect 29826 219200 29882 220000
rect 30838 219200 30894 220000
rect 31850 219200 31906 220000
rect 32862 219200 32918 220000
rect 33874 219200 33930 220000
rect 34886 219200 34942 220000
rect 35898 219200 35954 220000
rect 36910 219200 36966 220000
rect 37922 219200 37978 220000
rect 38934 219200 38990 220000
rect 39946 219200 40002 220000
rect 40958 219200 41014 220000
rect 41970 219200 42026 220000
rect 42982 219200 43038 220000
rect 43994 219200 44050 220000
rect 45006 219200 45062 220000
rect 46018 219200 46074 220000
rect 47030 219200 47086 220000
rect 48042 219200 48098 220000
rect 49054 219200 49110 220000
rect 50066 219200 50122 220000
rect 51078 219200 51134 220000
rect 52090 219200 52146 220000
rect 53102 219200 53158 220000
rect 54114 219200 54170 220000
rect 55126 219200 55182 220000
rect 56230 219200 56286 220000
rect 57242 219200 57298 220000
rect 58254 219200 58310 220000
rect 59266 219200 59322 220000
rect 60278 219200 60334 220000
rect 61290 219200 61346 220000
rect 62302 219200 62358 220000
rect 63314 219200 63370 220000
rect 64326 219200 64382 220000
rect 65338 219200 65394 220000
rect 66350 219200 66406 220000
rect 67362 219200 67418 220000
rect 68374 219200 68430 220000
rect 69386 219200 69442 220000
rect 70398 219200 70454 220000
rect 71410 219200 71466 220000
rect 72422 219200 72478 220000
rect 73434 219200 73490 220000
rect 74446 219200 74502 220000
rect 75458 219200 75514 220000
rect 76470 219200 76526 220000
rect 77482 219200 77538 220000
rect 78494 219200 78550 220000
rect 79506 219200 79562 220000
rect 80518 219200 80574 220000
rect 81530 219200 81586 220000
rect 82542 219200 82598 220000
rect 83554 219200 83610 220000
rect 84566 219200 84622 220000
rect 85578 219200 85634 220000
rect 86590 219200 86646 220000
rect 87602 219200 87658 220000
rect 88614 219200 88670 220000
rect 89626 219200 89682 220000
rect 90638 219200 90694 220000
rect 91650 219200 91706 220000
rect 92662 219200 92718 220000
rect 93674 219200 93730 220000
rect 94686 219200 94742 220000
rect 95698 219200 95754 220000
rect 96710 219200 96766 220000
rect 97722 219200 97778 220000
rect 98734 219200 98790 220000
rect 99746 219200 99802 220000
rect 100758 219200 100814 220000
rect 101770 219200 101826 220000
rect 102782 219200 102838 220000
rect 103794 219200 103850 220000
rect 104806 219200 104862 220000
rect 105818 219200 105874 220000
rect 106830 219200 106886 220000
rect 107842 219200 107898 220000
rect 108854 219200 108910 220000
rect 109866 219200 109922 220000
rect 110970 219200 111026 220000
rect 111982 219200 112038 220000
rect 112994 219200 113050 220000
rect 114006 219200 114062 220000
rect 115018 219200 115074 220000
rect 116030 219200 116086 220000
rect 117042 219200 117098 220000
rect 118054 219200 118110 220000
rect 119066 219200 119122 220000
rect 120078 219200 120134 220000
rect 121090 219200 121146 220000
rect 122102 219200 122158 220000
rect 123114 219200 123170 220000
rect 124126 219200 124182 220000
rect 125138 219200 125194 220000
rect 126150 219200 126206 220000
rect 127162 219200 127218 220000
rect 128174 219200 128230 220000
rect 129186 219200 129242 220000
rect 130198 219200 130254 220000
rect 131210 219200 131266 220000
rect 132222 219200 132278 220000
rect 133234 219200 133290 220000
rect 134246 219200 134302 220000
rect 135258 219200 135314 220000
rect 136270 219200 136326 220000
rect 137282 219200 137338 220000
rect 138294 219200 138350 220000
rect 139306 219200 139362 220000
rect 140318 219200 140374 220000
rect 141330 219200 141386 220000
rect 142342 219200 142398 220000
rect 143354 219200 143410 220000
rect 144366 219200 144422 220000
rect 145378 219200 145434 220000
rect 146390 219200 146446 220000
rect 147402 219200 147458 220000
rect 148414 219200 148470 220000
rect 149426 219200 149482 220000
rect 150438 219200 150494 220000
rect 151450 219200 151506 220000
rect 152462 219200 152518 220000
rect 153474 219200 153530 220000
rect 154486 219200 154542 220000
rect 155498 219200 155554 220000
rect 156510 219200 156566 220000
rect 157522 219200 157578 220000
rect 158534 219200 158590 220000
rect 159546 219200 159602 220000
rect 160558 219200 160614 220000
rect 161570 219200 161626 220000
rect 162582 219200 162638 220000
rect 163594 219200 163650 220000
rect 164606 219200 164662 220000
rect 165710 219200 165766 220000
rect 166722 219200 166778 220000
rect 167734 219200 167790 220000
rect 168746 219200 168802 220000
rect 169758 219200 169814 220000
rect 170770 219200 170826 220000
rect 171782 219200 171838 220000
rect 172794 219200 172850 220000
rect 173806 219200 173862 220000
rect 174818 219200 174874 220000
rect 175830 219200 175886 220000
rect 176842 219200 176898 220000
rect 177854 219200 177910 220000
rect 178866 219200 178922 220000
rect 179878 219200 179934 220000
rect 180890 219200 180946 220000
rect 181902 219200 181958 220000
rect 182914 219200 182970 220000
rect 183926 219200 183982 220000
rect 184938 219200 184994 220000
rect 185950 219200 186006 220000
rect 186962 219200 187018 220000
rect 187974 219200 188030 220000
rect 188986 219200 189042 220000
rect 189998 219200 190054 220000
rect 191010 219200 191066 220000
rect 192022 219200 192078 220000
rect 193034 219200 193090 220000
rect 194046 219200 194102 220000
rect 195058 219200 195114 220000
rect 196070 219200 196126 220000
rect 197082 219200 197138 220000
rect 198094 219200 198150 220000
rect 199106 219200 199162 220000
rect 200118 219200 200174 220000
rect 201130 219200 201186 220000
rect 202142 219200 202198 220000
rect 203154 219200 203210 220000
rect 204166 219200 204222 220000
rect 205178 219200 205234 220000
rect 206190 219200 206246 220000
rect 207202 219200 207258 220000
rect 208214 219200 208270 220000
rect 209226 219200 209282 220000
rect 210238 219200 210294 220000
rect 211250 219200 211306 220000
rect 212262 219200 212318 220000
rect 213274 219200 213330 220000
rect 214286 219200 214342 220000
rect 215298 219200 215354 220000
rect 216310 219200 216366 220000
rect 217322 219200 217378 220000
rect 218334 219200 218390 220000
rect 219346 219200 219402 220000
<< obsm2 >>
rect 18 219144 422 219200
rect 590 219144 1434 219200
rect 1602 219144 2446 219200
rect 2614 219144 3458 219200
rect 3626 219144 4470 219200
rect 4638 219144 5482 219200
rect 5650 219144 6494 219200
rect 6662 219144 7506 219200
rect 7674 219144 8518 219200
rect 8686 219144 9530 219200
rect 9698 219144 10542 219200
rect 10710 219144 11554 219200
rect 11722 219144 12566 219200
rect 12734 219144 13578 219200
rect 13746 219144 14590 219200
rect 14758 219144 15602 219200
rect 15770 219144 16614 219200
rect 16782 219144 17626 219200
rect 17794 219144 18638 219200
rect 18806 219144 19650 219200
rect 19818 219144 20662 219200
rect 20830 219144 21674 219200
rect 21842 219144 22686 219200
rect 22854 219144 23698 219200
rect 23866 219144 24710 219200
rect 24878 219144 25722 219200
rect 25890 219144 26734 219200
rect 26902 219144 27746 219200
rect 27914 219144 28758 219200
rect 28926 219144 29770 219200
rect 29938 219144 30782 219200
rect 30950 219144 31794 219200
rect 31962 219144 32806 219200
rect 32974 219144 33818 219200
rect 33986 219144 34830 219200
rect 34998 219144 35842 219200
rect 36010 219144 36854 219200
rect 37022 219144 37866 219200
rect 38034 219144 38878 219200
rect 39046 219144 39890 219200
rect 40058 219144 40902 219200
rect 41070 219144 41914 219200
rect 42082 219144 42926 219200
rect 43094 219144 43938 219200
rect 44106 219144 44950 219200
rect 45118 219144 45962 219200
rect 46130 219144 46974 219200
rect 47142 219144 47986 219200
rect 48154 219144 48998 219200
rect 49166 219144 50010 219200
rect 50178 219144 51022 219200
rect 51190 219144 52034 219200
rect 52202 219144 53046 219200
rect 53214 219144 54058 219200
rect 54226 219144 55070 219200
rect 55238 219144 56174 219200
rect 56342 219144 57186 219200
rect 57354 219144 58198 219200
rect 58366 219144 59210 219200
rect 59378 219144 60222 219200
rect 60390 219144 61234 219200
rect 61402 219144 62246 219200
rect 62414 219144 63258 219200
rect 63426 219144 64270 219200
rect 64438 219144 65282 219200
rect 65450 219144 66294 219200
rect 66462 219144 67306 219200
rect 67474 219144 68318 219200
rect 68486 219144 69330 219200
rect 69498 219144 70342 219200
rect 70510 219144 71354 219200
rect 71522 219144 72366 219200
rect 72534 219144 73378 219200
rect 73546 219144 74390 219200
rect 74558 219144 75402 219200
rect 75570 219144 76414 219200
rect 76582 219144 77426 219200
rect 77594 219144 78438 219200
rect 78606 219144 79450 219200
rect 79618 219144 80462 219200
rect 80630 219144 81474 219200
rect 81642 219144 82486 219200
rect 82654 219144 83498 219200
rect 83666 219144 84510 219200
rect 84678 219144 85522 219200
rect 85690 219144 86534 219200
rect 86702 219144 87546 219200
rect 87714 219144 88558 219200
rect 88726 219144 89570 219200
rect 89738 219144 90582 219200
rect 90750 219144 91594 219200
rect 91762 219144 92606 219200
rect 92774 219144 93618 219200
rect 93786 219144 94630 219200
rect 94798 219144 95642 219200
rect 95810 219144 96654 219200
rect 96822 219144 97666 219200
rect 97834 219144 98678 219200
rect 98846 219144 99690 219200
rect 99858 219144 100702 219200
rect 100870 219144 101714 219200
rect 101882 219144 102726 219200
rect 102894 219144 103738 219200
rect 103906 219144 104750 219200
rect 104918 219144 105762 219200
rect 105930 219144 106774 219200
rect 106942 219144 107786 219200
rect 107954 219144 108798 219200
rect 108966 219144 109810 219200
rect 109978 219144 110914 219200
rect 111082 219144 111926 219200
rect 112094 219144 112938 219200
rect 113106 219144 113950 219200
rect 114118 219144 114962 219200
rect 115130 219144 115974 219200
rect 116142 219144 116986 219200
rect 117154 219144 117998 219200
rect 118166 219144 119010 219200
rect 119178 219144 120022 219200
rect 120190 219144 121034 219200
rect 121202 219144 122046 219200
rect 122214 219144 123058 219200
rect 123226 219144 124070 219200
rect 124238 219144 125082 219200
rect 125250 219144 126094 219200
rect 126262 219144 127106 219200
rect 127274 219144 128118 219200
rect 128286 219144 129130 219200
rect 129298 219144 130142 219200
rect 130310 219144 131154 219200
rect 131322 219144 132166 219200
rect 132334 219144 133178 219200
rect 133346 219144 134190 219200
rect 134358 219144 135202 219200
rect 135370 219144 136214 219200
rect 136382 219144 137226 219200
rect 137394 219144 138238 219200
rect 138406 219144 139250 219200
rect 139418 219144 140262 219200
rect 140430 219144 141274 219200
rect 141442 219144 142286 219200
rect 142454 219144 143298 219200
rect 143466 219144 144310 219200
rect 144478 219144 145322 219200
rect 145490 219144 146334 219200
rect 146502 219144 147346 219200
rect 147514 219144 148358 219200
rect 148526 219144 149370 219200
rect 149538 219144 150382 219200
rect 150550 219144 151394 219200
rect 151562 219144 152406 219200
rect 152574 219144 153418 219200
rect 153586 219144 154430 219200
rect 154598 219144 155442 219200
rect 155610 219144 156454 219200
rect 156622 219144 157466 219200
rect 157634 219144 158478 219200
rect 158646 219144 159490 219200
rect 159658 219144 160502 219200
rect 160670 219144 161514 219200
rect 161682 219144 162526 219200
rect 162694 219144 163538 219200
rect 163706 219144 164550 219200
rect 164718 219144 165654 219200
rect 165822 219144 166666 219200
rect 166834 219144 167678 219200
rect 167846 219144 168690 219200
rect 168858 219144 169702 219200
rect 169870 219144 170714 219200
rect 170882 219144 171726 219200
rect 171894 219144 172738 219200
rect 172906 219144 173750 219200
rect 173918 219144 174762 219200
rect 174930 219144 175774 219200
rect 175942 219144 176786 219200
rect 176954 219144 177798 219200
rect 177966 219144 178810 219200
rect 178978 219144 179822 219200
rect 179990 219144 180834 219200
rect 181002 219144 181846 219200
rect 182014 219144 182858 219200
rect 183026 219144 183870 219200
rect 184038 219144 184882 219200
rect 185050 219144 185894 219200
rect 186062 219144 186906 219200
rect 187074 219144 187918 219200
rect 188086 219144 188930 219200
rect 189098 219144 189942 219200
rect 190110 219144 190954 219200
rect 191122 219144 191966 219200
rect 192134 219144 192978 219200
rect 193146 219144 193990 219200
rect 194158 219144 195002 219200
rect 195170 219144 196014 219200
rect 196182 219144 197026 219200
rect 197194 219144 198038 219200
rect 198206 219144 199050 219200
rect 199218 219144 200062 219200
rect 200230 219144 201074 219200
rect 201242 219144 202086 219200
rect 202254 219144 203098 219200
rect 203266 219144 204110 219200
rect 204278 219144 205122 219200
rect 205290 219144 206134 219200
rect 206302 219144 207146 219200
rect 207314 219144 208158 219200
rect 208326 219144 209170 219200
rect 209338 219144 210182 219200
rect 210350 219144 211194 219200
rect 211362 219144 212206 219200
rect 212374 219144 213218 219200
rect 213386 219144 214230 219200
rect 214398 219144 215242 219200
rect 215410 219144 216254 219200
rect 216422 219144 217266 219200
rect 217434 219144 218278 219200
rect 218446 219144 219290 219200
rect 18 2128 219400 219144
<< metal3 >>
rect 0 218424 800 218544
rect 0 215432 800 215552
rect 0 212304 800 212424
rect 0 209312 800 209432
rect 0 206184 800 206304
rect 0 203192 800 203312
rect 0 200064 800 200184
rect 0 197072 800 197192
rect 0 193944 800 194064
rect 0 190952 800 191072
rect 0 187824 800 187944
rect 0 184832 800 184952
rect 0 181704 800 181824
rect 0 178712 800 178832
rect 0 175584 800 175704
rect 0 172592 800 172712
rect 0 169464 800 169584
rect 0 166472 800 166592
rect 0 163480 800 163600
rect 0 160352 800 160472
rect 0 157360 800 157480
rect 0 154232 800 154352
rect 0 151240 800 151360
rect 0 148112 800 148232
rect 0 145120 800 145240
rect 0 141992 800 142112
rect 0 139000 800 139120
rect 0 135872 800 135992
rect 0 132880 800 133000
rect 0 129752 800 129872
rect 0 126760 800 126880
rect 0 123632 800 123752
rect 0 120640 800 120760
rect 0 117512 800 117632
rect 0 114520 800 114640
rect 0 111528 800 111648
rect 0 108400 800 108520
rect 0 105408 800 105528
rect 0 102280 800 102400
rect 0 99288 800 99408
rect 0 96160 800 96280
rect 0 93168 800 93288
rect 0 90040 800 90160
rect 0 87048 800 87168
rect 0 83920 800 84040
rect 0 80928 800 81048
rect 0 77800 800 77920
rect 0 74808 800 74928
rect 0 71680 800 71800
rect 0 68688 800 68808
rect 0 65560 800 65680
rect 0 62568 800 62688
rect 0 59440 800 59560
rect 0 56448 800 56568
rect 0 53456 800 53576
rect 0 50328 800 50448
rect 0 47336 800 47456
rect 0 44208 800 44328
rect 0 41216 800 41336
rect 0 38088 800 38208
rect 0 35096 800 35216
rect 0 31968 800 32088
rect 0 28976 800 29096
rect 0 25848 800 25968
rect 0 22856 800 22976
rect 0 19728 800 19848
rect 0 16736 800 16856
rect 0 13608 800 13728
rect 0 10616 800 10736
rect 0 7488 800 7608
rect 0 4496 800 4616
rect 0 1504 800 1624
<< obsm3 >>
rect 880 218344 218487 218514
rect 13 215632 218487 218344
rect 880 215352 218487 215632
rect 13 212504 218487 215352
rect 880 212224 218487 212504
rect 13 209512 218487 212224
rect 880 209232 218487 209512
rect 13 206384 218487 209232
rect 880 206104 218487 206384
rect 13 203392 218487 206104
rect 880 203112 218487 203392
rect 13 200264 218487 203112
rect 880 199984 218487 200264
rect 13 197272 218487 199984
rect 880 196992 218487 197272
rect 13 194144 218487 196992
rect 880 193864 218487 194144
rect 13 191152 218487 193864
rect 880 190872 218487 191152
rect 13 188024 218487 190872
rect 880 187744 218487 188024
rect 13 185032 218487 187744
rect 880 184752 218487 185032
rect 13 181904 218487 184752
rect 880 181624 218487 181904
rect 13 178912 218487 181624
rect 880 178632 218487 178912
rect 13 175784 218487 178632
rect 880 175504 218487 175784
rect 13 172792 218487 175504
rect 880 172512 218487 172792
rect 13 169664 218487 172512
rect 880 169384 218487 169664
rect 13 166672 218487 169384
rect 880 166392 218487 166672
rect 13 163680 218487 166392
rect 880 163400 218487 163680
rect 13 160552 218487 163400
rect 880 160272 218487 160552
rect 13 157560 218487 160272
rect 880 157280 218487 157560
rect 13 154432 218487 157280
rect 880 154152 218487 154432
rect 13 151440 218487 154152
rect 880 151160 218487 151440
rect 13 148312 218487 151160
rect 880 148032 218487 148312
rect 13 145320 218487 148032
rect 880 145040 218487 145320
rect 13 142192 218487 145040
rect 880 141912 218487 142192
rect 13 139200 218487 141912
rect 880 138920 218487 139200
rect 13 136072 218487 138920
rect 880 135792 218487 136072
rect 13 133080 218487 135792
rect 880 132800 218487 133080
rect 13 129952 218487 132800
rect 880 129672 218487 129952
rect 13 126960 218487 129672
rect 880 126680 218487 126960
rect 13 123832 218487 126680
rect 880 123552 218487 123832
rect 13 120840 218487 123552
rect 880 120560 218487 120840
rect 13 117712 218487 120560
rect 880 117432 218487 117712
rect 13 114720 218487 117432
rect 880 114440 218487 114720
rect 13 111728 218487 114440
rect 880 111448 218487 111728
rect 13 108600 218487 111448
rect 880 108320 218487 108600
rect 13 105608 218487 108320
rect 880 105328 218487 105608
rect 13 102480 218487 105328
rect 880 102200 218487 102480
rect 13 99488 218487 102200
rect 880 99208 218487 99488
rect 13 96360 218487 99208
rect 880 96080 218487 96360
rect 13 93368 218487 96080
rect 880 93088 218487 93368
rect 13 90240 218487 93088
rect 880 89960 218487 90240
rect 13 87248 218487 89960
rect 880 86968 218487 87248
rect 13 84120 218487 86968
rect 880 83840 218487 84120
rect 13 81128 218487 83840
rect 880 80848 218487 81128
rect 13 78000 218487 80848
rect 880 77720 218487 78000
rect 13 75008 218487 77720
rect 880 74728 218487 75008
rect 13 71880 218487 74728
rect 880 71600 218487 71880
rect 13 68888 218487 71600
rect 880 68608 218487 68888
rect 13 65760 218487 68608
rect 880 65480 218487 65760
rect 13 62768 218487 65480
rect 880 62488 218487 62768
rect 13 59640 218487 62488
rect 880 59360 218487 59640
rect 13 56648 218487 59360
rect 880 56368 218487 56648
rect 13 53656 218487 56368
rect 880 53376 218487 53656
rect 13 50528 218487 53376
rect 880 50248 218487 50528
rect 13 47536 218487 50248
rect 880 47256 218487 47536
rect 13 44408 218487 47256
rect 880 44128 218487 44408
rect 13 41416 218487 44128
rect 880 41136 218487 41416
rect 13 38288 218487 41136
rect 880 38008 218487 38288
rect 13 35296 218487 38008
rect 880 35016 218487 35296
rect 13 32168 218487 35016
rect 880 31888 218487 32168
rect 13 29176 218487 31888
rect 880 28896 218487 29176
rect 13 26048 218487 28896
rect 880 25768 218487 26048
rect 13 23056 218487 25768
rect 880 22776 218487 23056
rect 13 19928 218487 22776
rect 880 19648 218487 19928
rect 13 16936 218487 19648
rect 880 16656 218487 16936
rect 13 13808 218487 16656
rect 880 13528 218487 13808
rect 13 10816 218487 13528
rect 880 10536 218487 10816
rect 13 7688 218487 10536
rect 880 7408 218487 7688
rect 13 4696 218487 7408
rect 880 4416 218487 4696
rect 13 1704 218487 4416
rect 880 1532 218487 1704
<< metal4 >>
rect 4208 2128 4528 217648
rect 19568 2128 19888 217648
rect 34928 2128 35248 217648
rect 50288 2128 50608 217648
rect 65648 2128 65968 217648
rect 81008 2128 81328 217648
rect 96368 2128 96688 217648
rect 111728 2128 112048 217648
rect 127088 2128 127408 217648
rect 142448 2128 142768 217648
rect 157808 2128 158128 217648
rect 173168 2128 173488 217648
rect 188528 2128 188848 217648
rect 203888 2128 204208 217648
<< obsm4 >>
rect 1715 217728 217797 217973
rect 1715 2048 4128 217728
rect 4608 2048 19488 217728
rect 19968 2048 34848 217728
rect 35328 2048 50208 217728
rect 50688 2048 65568 217728
rect 66048 2048 80928 217728
rect 81408 2048 96288 217728
rect 96768 2048 111648 217728
rect 112128 2048 127008 217728
rect 127488 2048 142368 217728
rect 142848 2048 157728 217728
rect 158208 2048 173088 217728
rect 173568 2048 188448 217728
rect 188928 2048 203808 217728
rect 204288 2048 217797 217728
rect 1715 1531 217797 2048
<< labels >>
rlabel metal2 s 478 219200 534 220000 6 clk
port 1 nsew signal input
rlabel metal2 s 1490 219200 1546 220000 6 d_in[0]
port 2 nsew signal input
rlabel metal2 s 11610 219200 11666 220000 6 d_in[10]
port 3 nsew signal input
rlabel metal2 s 12622 219200 12678 220000 6 d_in[11]
port 4 nsew signal input
rlabel metal2 s 13634 219200 13690 220000 6 d_in[12]
port 5 nsew signal input
rlabel metal2 s 14646 219200 14702 220000 6 d_in[13]
port 6 nsew signal input
rlabel metal2 s 15658 219200 15714 220000 6 d_in[14]
port 7 nsew signal input
rlabel metal2 s 16670 219200 16726 220000 6 d_in[15]
port 8 nsew signal input
rlabel metal2 s 17682 219200 17738 220000 6 d_in[16]
port 9 nsew signal input
rlabel metal2 s 18694 219200 18750 220000 6 d_in[17]
port 10 nsew signal input
rlabel metal2 s 19706 219200 19762 220000 6 d_in[18]
port 11 nsew signal input
rlabel metal2 s 20718 219200 20774 220000 6 d_in[19]
port 12 nsew signal input
rlabel metal2 s 2502 219200 2558 220000 6 d_in[1]
port 13 nsew signal input
rlabel metal2 s 21730 219200 21786 220000 6 d_in[20]
port 14 nsew signal input
rlabel metal2 s 22742 219200 22798 220000 6 d_in[21]
port 15 nsew signal input
rlabel metal2 s 23754 219200 23810 220000 6 d_in[22]
port 16 nsew signal input
rlabel metal2 s 24766 219200 24822 220000 6 d_in[23]
port 17 nsew signal input
rlabel metal2 s 3514 219200 3570 220000 6 d_in[2]
port 18 nsew signal input
rlabel metal2 s 4526 219200 4582 220000 6 d_in[3]
port 19 nsew signal input
rlabel metal2 s 5538 219200 5594 220000 6 d_in[4]
port 20 nsew signal input
rlabel metal2 s 6550 219200 6606 220000 6 d_in[5]
port 21 nsew signal input
rlabel metal2 s 7562 219200 7618 220000 6 d_in[6]
port 22 nsew signal input
rlabel metal2 s 8574 219200 8630 220000 6 d_in[7]
port 23 nsew signal input
rlabel metal2 s 9586 219200 9642 220000 6 d_in[8]
port 24 nsew signal input
rlabel metal2 s 10598 219200 10654 220000 6 d_in[9]
port 25 nsew signal input
rlabel metal2 s 25778 219200 25834 220000 6 d_out[0]
port 26 nsew signal output
rlabel metal2 s 127162 219200 127218 220000 6 d_out[100]
port 27 nsew signal output
rlabel metal2 s 128174 219200 128230 220000 6 d_out[101]
port 28 nsew signal output
rlabel metal2 s 129186 219200 129242 220000 6 d_out[102]
port 29 nsew signal output
rlabel metal2 s 130198 219200 130254 220000 6 d_out[103]
port 30 nsew signal output
rlabel metal2 s 131210 219200 131266 220000 6 d_out[104]
port 31 nsew signal output
rlabel metal2 s 132222 219200 132278 220000 6 d_out[105]
port 32 nsew signal output
rlabel metal2 s 133234 219200 133290 220000 6 d_out[106]
port 33 nsew signal output
rlabel metal2 s 134246 219200 134302 220000 6 d_out[107]
port 34 nsew signal output
rlabel metal2 s 135258 219200 135314 220000 6 d_out[108]
port 35 nsew signal output
rlabel metal2 s 136270 219200 136326 220000 6 d_out[109]
port 36 nsew signal output
rlabel metal2 s 35898 219200 35954 220000 6 d_out[10]
port 37 nsew signal output
rlabel metal2 s 137282 219200 137338 220000 6 d_out[110]
port 38 nsew signal output
rlabel metal2 s 138294 219200 138350 220000 6 d_out[111]
port 39 nsew signal output
rlabel metal2 s 139306 219200 139362 220000 6 d_out[112]
port 40 nsew signal output
rlabel metal2 s 140318 219200 140374 220000 6 d_out[113]
port 41 nsew signal output
rlabel metal2 s 141330 219200 141386 220000 6 d_out[114]
port 42 nsew signal output
rlabel metal2 s 142342 219200 142398 220000 6 d_out[115]
port 43 nsew signal output
rlabel metal2 s 143354 219200 143410 220000 6 d_out[116]
port 44 nsew signal output
rlabel metal2 s 144366 219200 144422 220000 6 d_out[117]
port 45 nsew signal output
rlabel metal2 s 145378 219200 145434 220000 6 d_out[118]
port 46 nsew signal output
rlabel metal2 s 146390 219200 146446 220000 6 d_out[119]
port 47 nsew signal output
rlabel metal2 s 36910 219200 36966 220000 6 d_out[11]
port 48 nsew signal output
rlabel metal2 s 147402 219200 147458 220000 6 d_out[120]
port 49 nsew signal output
rlabel metal2 s 148414 219200 148470 220000 6 d_out[121]
port 50 nsew signal output
rlabel metal2 s 149426 219200 149482 220000 6 d_out[122]
port 51 nsew signal output
rlabel metal2 s 150438 219200 150494 220000 6 d_out[123]
port 52 nsew signal output
rlabel metal2 s 151450 219200 151506 220000 6 d_out[124]
port 53 nsew signal output
rlabel metal2 s 152462 219200 152518 220000 6 d_out[125]
port 54 nsew signal output
rlabel metal2 s 153474 219200 153530 220000 6 d_out[126]
port 55 nsew signal output
rlabel metal2 s 154486 219200 154542 220000 6 d_out[127]
port 56 nsew signal output
rlabel metal2 s 155498 219200 155554 220000 6 d_out[128]
port 57 nsew signal output
rlabel metal2 s 156510 219200 156566 220000 6 d_out[129]
port 58 nsew signal output
rlabel metal2 s 37922 219200 37978 220000 6 d_out[12]
port 59 nsew signal output
rlabel metal2 s 157522 219200 157578 220000 6 d_out[130]
port 60 nsew signal output
rlabel metal2 s 158534 219200 158590 220000 6 d_out[131]
port 61 nsew signal output
rlabel metal2 s 159546 219200 159602 220000 6 d_out[132]
port 62 nsew signal output
rlabel metal2 s 160558 219200 160614 220000 6 d_out[133]
port 63 nsew signal output
rlabel metal2 s 161570 219200 161626 220000 6 d_out[134]
port 64 nsew signal output
rlabel metal2 s 162582 219200 162638 220000 6 d_out[135]
port 65 nsew signal output
rlabel metal2 s 163594 219200 163650 220000 6 d_out[136]
port 66 nsew signal output
rlabel metal2 s 164606 219200 164662 220000 6 d_out[137]
port 67 nsew signal output
rlabel metal2 s 165710 219200 165766 220000 6 d_out[138]
port 68 nsew signal output
rlabel metal2 s 166722 219200 166778 220000 6 d_out[139]
port 69 nsew signal output
rlabel metal2 s 38934 219200 38990 220000 6 d_out[13]
port 70 nsew signal output
rlabel metal2 s 167734 219200 167790 220000 6 d_out[140]
port 71 nsew signal output
rlabel metal2 s 168746 219200 168802 220000 6 d_out[141]
port 72 nsew signal output
rlabel metal2 s 169758 219200 169814 220000 6 d_out[142]
port 73 nsew signal output
rlabel metal2 s 170770 219200 170826 220000 6 d_out[143]
port 74 nsew signal output
rlabel metal2 s 171782 219200 171838 220000 6 d_out[144]
port 75 nsew signal output
rlabel metal2 s 172794 219200 172850 220000 6 d_out[145]
port 76 nsew signal output
rlabel metal2 s 173806 219200 173862 220000 6 d_out[146]
port 77 nsew signal output
rlabel metal2 s 174818 219200 174874 220000 6 d_out[147]
port 78 nsew signal output
rlabel metal2 s 175830 219200 175886 220000 6 d_out[148]
port 79 nsew signal output
rlabel metal2 s 176842 219200 176898 220000 6 d_out[149]
port 80 nsew signal output
rlabel metal2 s 39946 219200 40002 220000 6 d_out[14]
port 81 nsew signal output
rlabel metal2 s 177854 219200 177910 220000 6 d_out[150]
port 82 nsew signal output
rlabel metal2 s 178866 219200 178922 220000 6 d_out[151]
port 83 nsew signal output
rlabel metal2 s 179878 219200 179934 220000 6 d_out[152]
port 84 nsew signal output
rlabel metal2 s 180890 219200 180946 220000 6 d_out[153]
port 85 nsew signal output
rlabel metal2 s 181902 219200 181958 220000 6 d_out[154]
port 86 nsew signal output
rlabel metal2 s 182914 219200 182970 220000 6 d_out[155]
port 87 nsew signal output
rlabel metal2 s 183926 219200 183982 220000 6 d_out[156]
port 88 nsew signal output
rlabel metal2 s 184938 219200 184994 220000 6 d_out[157]
port 89 nsew signal output
rlabel metal2 s 185950 219200 186006 220000 6 d_out[158]
port 90 nsew signal output
rlabel metal2 s 186962 219200 187018 220000 6 d_out[159]
port 91 nsew signal output
rlabel metal2 s 40958 219200 41014 220000 6 d_out[15]
port 92 nsew signal output
rlabel metal2 s 187974 219200 188030 220000 6 d_out[160]
port 93 nsew signal output
rlabel metal2 s 188986 219200 189042 220000 6 d_out[161]
port 94 nsew signal output
rlabel metal2 s 189998 219200 190054 220000 6 d_out[162]
port 95 nsew signal output
rlabel metal2 s 191010 219200 191066 220000 6 d_out[163]
port 96 nsew signal output
rlabel metal2 s 192022 219200 192078 220000 6 d_out[164]
port 97 nsew signal output
rlabel metal2 s 193034 219200 193090 220000 6 d_out[165]
port 98 nsew signal output
rlabel metal2 s 194046 219200 194102 220000 6 d_out[166]
port 99 nsew signal output
rlabel metal2 s 195058 219200 195114 220000 6 d_out[167]
port 100 nsew signal output
rlabel metal2 s 196070 219200 196126 220000 6 d_out[168]
port 101 nsew signal output
rlabel metal2 s 197082 219200 197138 220000 6 d_out[169]
port 102 nsew signal output
rlabel metal2 s 41970 219200 42026 220000 6 d_out[16]
port 103 nsew signal output
rlabel metal2 s 198094 219200 198150 220000 6 d_out[170]
port 104 nsew signal output
rlabel metal2 s 199106 219200 199162 220000 6 d_out[171]
port 105 nsew signal output
rlabel metal2 s 200118 219200 200174 220000 6 d_out[172]
port 106 nsew signal output
rlabel metal2 s 201130 219200 201186 220000 6 d_out[173]
port 107 nsew signal output
rlabel metal2 s 202142 219200 202198 220000 6 d_out[174]
port 108 nsew signal output
rlabel metal2 s 203154 219200 203210 220000 6 d_out[175]
port 109 nsew signal output
rlabel metal2 s 204166 219200 204222 220000 6 d_out[176]
port 110 nsew signal output
rlabel metal2 s 205178 219200 205234 220000 6 d_out[177]
port 111 nsew signal output
rlabel metal2 s 206190 219200 206246 220000 6 d_out[178]
port 112 nsew signal output
rlabel metal2 s 207202 219200 207258 220000 6 d_out[179]
port 113 nsew signal output
rlabel metal2 s 42982 219200 43038 220000 6 d_out[17]
port 114 nsew signal output
rlabel metal2 s 208214 219200 208270 220000 6 d_out[180]
port 115 nsew signal output
rlabel metal2 s 209226 219200 209282 220000 6 d_out[181]
port 116 nsew signal output
rlabel metal2 s 210238 219200 210294 220000 6 d_out[182]
port 117 nsew signal output
rlabel metal2 s 211250 219200 211306 220000 6 d_out[183]
port 118 nsew signal output
rlabel metal2 s 212262 219200 212318 220000 6 d_out[184]
port 119 nsew signal output
rlabel metal2 s 213274 219200 213330 220000 6 d_out[185]
port 120 nsew signal output
rlabel metal2 s 214286 219200 214342 220000 6 d_out[186]
port 121 nsew signal output
rlabel metal2 s 215298 219200 215354 220000 6 d_out[187]
port 122 nsew signal output
rlabel metal2 s 216310 219200 216366 220000 6 d_out[188]
port 123 nsew signal output
rlabel metal2 s 217322 219200 217378 220000 6 d_out[189]
port 124 nsew signal output
rlabel metal2 s 43994 219200 44050 220000 6 d_out[18]
port 125 nsew signal output
rlabel metal2 s 218334 219200 218390 220000 6 d_out[190]
port 126 nsew signal output
rlabel metal2 s 219346 219200 219402 220000 6 d_out[191]
port 127 nsew signal output
rlabel metal2 s 45006 219200 45062 220000 6 d_out[19]
port 128 nsew signal output
rlabel metal2 s 26790 219200 26846 220000 6 d_out[1]
port 129 nsew signal output
rlabel metal2 s 46018 219200 46074 220000 6 d_out[20]
port 130 nsew signal output
rlabel metal2 s 47030 219200 47086 220000 6 d_out[21]
port 131 nsew signal output
rlabel metal2 s 48042 219200 48098 220000 6 d_out[22]
port 132 nsew signal output
rlabel metal2 s 49054 219200 49110 220000 6 d_out[23]
port 133 nsew signal output
rlabel metal2 s 50066 219200 50122 220000 6 d_out[24]
port 134 nsew signal output
rlabel metal2 s 51078 219200 51134 220000 6 d_out[25]
port 135 nsew signal output
rlabel metal2 s 52090 219200 52146 220000 6 d_out[26]
port 136 nsew signal output
rlabel metal2 s 53102 219200 53158 220000 6 d_out[27]
port 137 nsew signal output
rlabel metal2 s 54114 219200 54170 220000 6 d_out[28]
port 138 nsew signal output
rlabel metal2 s 55126 219200 55182 220000 6 d_out[29]
port 139 nsew signal output
rlabel metal2 s 27802 219200 27858 220000 6 d_out[2]
port 140 nsew signal output
rlabel metal2 s 56230 219200 56286 220000 6 d_out[30]
port 141 nsew signal output
rlabel metal2 s 57242 219200 57298 220000 6 d_out[31]
port 142 nsew signal output
rlabel metal2 s 58254 219200 58310 220000 6 d_out[32]
port 143 nsew signal output
rlabel metal2 s 59266 219200 59322 220000 6 d_out[33]
port 144 nsew signal output
rlabel metal2 s 60278 219200 60334 220000 6 d_out[34]
port 145 nsew signal output
rlabel metal2 s 61290 219200 61346 220000 6 d_out[35]
port 146 nsew signal output
rlabel metal2 s 62302 219200 62358 220000 6 d_out[36]
port 147 nsew signal output
rlabel metal2 s 63314 219200 63370 220000 6 d_out[37]
port 148 nsew signal output
rlabel metal2 s 64326 219200 64382 220000 6 d_out[38]
port 149 nsew signal output
rlabel metal2 s 65338 219200 65394 220000 6 d_out[39]
port 150 nsew signal output
rlabel metal2 s 28814 219200 28870 220000 6 d_out[3]
port 151 nsew signal output
rlabel metal2 s 66350 219200 66406 220000 6 d_out[40]
port 152 nsew signal output
rlabel metal2 s 67362 219200 67418 220000 6 d_out[41]
port 153 nsew signal output
rlabel metal2 s 68374 219200 68430 220000 6 d_out[42]
port 154 nsew signal output
rlabel metal2 s 69386 219200 69442 220000 6 d_out[43]
port 155 nsew signal output
rlabel metal2 s 70398 219200 70454 220000 6 d_out[44]
port 156 nsew signal output
rlabel metal2 s 71410 219200 71466 220000 6 d_out[45]
port 157 nsew signal output
rlabel metal2 s 72422 219200 72478 220000 6 d_out[46]
port 158 nsew signal output
rlabel metal2 s 73434 219200 73490 220000 6 d_out[47]
port 159 nsew signal output
rlabel metal2 s 74446 219200 74502 220000 6 d_out[48]
port 160 nsew signal output
rlabel metal2 s 75458 219200 75514 220000 6 d_out[49]
port 161 nsew signal output
rlabel metal2 s 29826 219200 29882 220000 6 d_out[4]
port 162 nsew signal output
rlabel metal2 s 76470 219200 76526 220000 6 d_out[50]
port 163 nsew signal output
rlabel metal2 s 77482 219200 77538 220000 6 d_out[51]
port 164 nsew signal output
rlabel metal2 s 78494 219200 78550 220000 6 d_out[52]
port 165 nsew signal output
rlabel metal2 s 79506 219200 79562 220000 6 d_out[53]
port 166 nsew signal output
rlabel metal2 s 80518 219200 80574 220000 6 d_out[54]
port 167 nsew signal output
rlabel metal2 s 81530 219200 81586 220000 6 d_out[55]
port 168 nsew signal output
rlabel metal2 s 82542 219200 82598 220000 6 d_out[56]
port 169 nsew signal output
rlabel metal2 s 83554 219200 83610 220000 6 d_out[57]
port 170 nsew signal output
rlabel metal2 s 84566 219200 84622 220000 6 d_out[58]
port 171 nsew signal output
rlabel metal2 s 85578 219200 85634 220000 6 d_out[59]
port 172 nsew signal output
rlabel metal2 s 30838 219200 30894 220000 6 d_out[5]
port 173 nsew signal output
rlabel metal2 s 86590 219200 86646 220000 6 d_out[60]
port 174 nsew signal output
rlabel metal2 s 87602 219200 87658 220000 6 d_out[61]
port 175 nsew signal output
rlabel metal2 s 88614 219200 88670 220000 6 d_out[62]
port 176 nsew signal output
rlabel metal2 s 89626 219200 89682 220000 6 d_out[63]
port 177 nsew signal output
rlabel metal2 s 90638 219200 90694 220000 6 d_out[64]
port 178 nsew signal output
rlabel metal2 s 91650 219200 91706 220000 6 d_out[65]
port 179 nsew signal output
rlabel metal2 s 92662 219200 92718 220000 6 d_out[66]
port 180 nsew signal output
rlabel metal2 s 93674 219200 93730 220000 6 d_out[67]
port 181 nsew signal output
rlabel metal2 s 94686 219200 94742 220000 6 d_out[68]
port 182 nsew signal output
rlabel metal2 s 95698 219200 95754 220000 6 d_out[69]
port 183 nsew signal output
rlabel metal2 s 31850 219200 31906 220000 6 d_out[6]
port 184 nsew signal output
rlabel metal2 s 96710 219200 96766 220000 6 d_out[70]
port 185 nsew signal output
rlabel metal2 s 97722 219200 97778 220000 6 d_out[71]
port 186 nsew signal output
rlabel metal2 s 98734 219200 98790 220000 6 d_out[72]
port 187 nsew signal output
rlabel metal2 s 99746 219200 99802 220000 6 d_out[73]
port 188 nsew signal output
rlabel metal2 s 100758 219200 100814 220000 6 d_out[74]
port 189 nsew signal output
rlabel metal2 s 101770 219200 101826 220000 6 d_out[75]
port 190 nsew signal output
rlabel metal2 s 102782 219200 102838 220000 6 d_out[76]
port 191 nsew signal output
rlabel metal2 s 103794 219200 103850 220000 6 d_out[77]
port 192 nsew signal output
rlabel metal2 s 104806 219200 104862 220000 6 d_out[78]
port 193 nsew signal output
rlabel metal2 s 105818 219200 105874 220000 6 d_out[79]
port 194 nsew signal output
rlabel metal2 s 32862 219200 32918 220000 6 d_out[7]
port 195 nsew signal output
rlabel metal2 s 106830 219200 106886 220000 6 d_out[80]
port 196 nsew signal output
rlabel metal2 s 107842 219200 107898 220000 6 d_out[81]
port 197 nsew signal output
rlabel metal2 s 108854 219200 108910 220000 6 d_out[82]
port 198 nsew signal output
rlabel metal2 s 109866 219200 109922 220000 6 d_out[83]
port 199 nsew signal output
rlabel metal2 s 110970 219200 111026 220000 6 d_out[84]
port 200 nsew signal output
rlabel metal2 s 111982 219200 112038 220000 6 d_out[85]
port 201 nsew signal output
rlabel metal2 s 112994 219200 113050 220000 6 d_out[86]
port 202 nsew signal output
rlabel metal2 s 114006 219200 114062 220000 6 d_out[87]
port 203 nsew signal output
rlabel metal2 s 115018 219200 115074 220000 6 d_out[88]
port 204 nsew signal output
rlabel metal2 s 116030 219200 116086 220000 6 d_out[89]
port 205 nsew signal output
rlabel metal2 s 33874 219200 33930 220000 6 d_out[8]
port 206 nsew signal output
rlabel metal2 s 117042 219200 117098 220000 6 d_out[90]
port 207 nsew signal output
rlabel metal2 s 118054 219200 118110 220000 6 d_out[91]
port 208 nsew signal output
rlabel metal2 s 119066 219200 119122 220000 6 d_out[92]
port 209 nsew signal output
rlabel metal2 s 120078 219200 120134 220000 6 d_out[93]
port 210 nsew signal output
rlabel metal2 s 121090 219200 121146 220000 6 d_out[94]
port 211 nsew signal output
rlabel metal2 s 122102 219200 122158 220000 6 d_out[95]
port 212 nsew signal output
rlabel metal2 s 123114 219200 123170 220000 6 d_out[96]
port 213 nsew signal output
rlabel metal2 s 124126 219200 124182 220000 6 d_out[97]
port 214 nsew signal output
rlabel metal2 s 125138 219200 125194 220000 6 d_out[98]
port 215 nsew signal output
rlabel metal2 s 126150 219200 126206 220000 6 d_out[99]
port 216 nsew signal output
rlabel metal2 s 34886 219200 34942 220000 6 d_out[9]
port 217 nsew signal output
rlabel metal3 s 0 1504 800 1624 6 w_in[0]
port 218 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 w_in[10]
port 219 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 w_in[11]
port 220 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 w_in[12]
port 221 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 w_in[13]
port 222 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 w_in[14]
port 223 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 w_in[15]
port 224 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 w_in[16]
port 225 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 w_in[17]
port 226 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 w_in[18]
port 227 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 w_in[19]
port 228 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 w_in[1]
port 229 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 w_in[20]
port 230 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 w_in[21]
port 231 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 w_in[22]
port 232 nsew signal input
rlabel metal3 s 0 71680 800 71800 6 w_in[23]
port 233 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 w_in[24]
port 234 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 w_in[25]
port 235 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 w_in[26]
port 236 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 w_in[27]
port 237 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 w_in[28]
port 238 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 w_in[29]
port 239 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 w_in[2]
port 240 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 w_in[30]
port 241 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 w_in[31]
port 242 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 w_in[32]
port 243 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 w_in[33]
port 244 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 w_in[34]
port 245 nsew signal input
rlabel metal3 s 0 108400 800 108520 6 w_in[35]
port 246 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 w_in[36]
port 247 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 w_in[37]
port 248 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 w_in[38]
port 249 nsew signal input
rlabel metal3 s 0 120640 800 120760 6 w_in[39]
port 250 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 w_in[3]
port 251 nsew signal input
rlabel metal3 s 0 123632 800 123752 6 w_in[40]
port 252 nsew signal input
rlabel metal3 s 0 126760 800 126880 6 w_in[41]
port 253 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 w_in[42]
port 254 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 w_in[43]
port 255 nsew signal input
rlabel metal3 s 0 135872 800 135992 6 w_in[44]
port 256 nsew signal input
rlabel metal3 s 0 139000 800 139120 6 w_in[45]
port 257 nsew signal input
rlabel metal3 s 0 141992 800 142112 6 w_in[46]
port 258 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 w_in[47]
port 259 nsew signal input
rlabel metal3 s 0 148112 800 148232 6 w_in[48]
port 260 nsew signal input
rlabel metal3 s 0 151240 800 151360 6 w_in[49]
port 261 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 w_in[4]
port 262 nsew signal input
rlabel metal3 s 0 154232 800 154352 6 w_in[50]
port 263 nsew signal input
rlabel metal3 s 0 157360 800 157480 6 w_in[51]
port 264 nsew signal input
rlabel metal3 s 0 160352 800 160472 6 w_in[52]
port 265 nsew signal input
rlabel metal3 s 0 163480 800 163600 6 w_in[53]
port 266 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 w_in[54]
port 267 nsew signal input
rlabel metal3 s 0 169464 800 169584 6 w_in[55]
port 268 nsew signal input
rlabel metal3 s 0 172592 800 172712 6 w_in[56]
port 269 nsew signal input
rlabel metal3 s 0 175584 800 175704 6 w_in[57]
port 270 nsew signal input
rlabel metal3 s 0 178712 800 178832 6 w_in[58]
port 271 nsew signal input
rlabel metal3 s 0 181704 800 181824 6 w_in[59]
port 272 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 w_in[5]
port 273 nsew signal input
rlabel metal3 s 0 184832 800 184952 6 w_in[60]
port 274 nsew signal input
rlabel metal3 s 0 187824 800 187944 6 w_in[61]
port 275 nsew signal input
rlabel metal3 s 0 190952 800 191072 6 w_in[62]
port 276 nsew signal input
rlabel metal3 s 0 193944 800 194064 6 w_in[63]
port 277 nsew signal input
rlabel metal3 s 0 197072 800 197192 6 w_in[64]
port 278 nsew signal input
rlabel metal3 s 0 200064 800 200184 6 w_in[65]
port 279 nsew signal input
rlabel metal3 s 0 203192 800 203312 6 w_in[66]
port 280 nsew signal input
rlabel metal3 s 0 206184 800 206304 6 w_in[67]
port 281 nsew signal input
rlabel metal3 s 0 209312 800 209432 6 w_in[68]
port 282 nsew signal input
rlabel metal3 s 0 212304 800 212424 6 w_in[69]
port 283 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 w_in[6]
port 284 nsew signal input
rlabel metal3 s 0 215432 800 215552 6 w_in[70]
port 285 nsew signal input
rlabel metal3 s 0 218424 800 218544 6 w_in[71]
port 286 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 w_in[7]
port 287 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 w_in[8]
port 288 nsew signal input
rlabel metal3 s 0 28976 800 29096 6 w_in[9]
port 289 nsew signal input
rlabel metal4 s 188528 2128 188848 217648 6 vccd1
port 290 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 217648 6 vccd1
port 291 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 217648 6 vccd1
port 292 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 217648 6 vccd1
port 293 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 217648 6 vccd1
port 294 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 217648 6 vccd1
port 295 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 217648 6 vccd1
port 296 nsew power bidirectional
rlabel metal4 s 203888 2128 204208 217648 6 vssd1
port 297 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 217648 6 vssd1
port 298 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 217648 6 vssd1
port 299 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 217648 6 vssd1
port 300 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 217648 6 vssd1
port 301 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 217648 6 vssd1
port 302 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 217648 6 vssd1
port 303 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 220000 220000
string LEFview TRUE
string GDS_FILE /project/openlane/register_file/runs/register_file/results/magic/register_file.gds
string GDS_END 151935626
string GDS_START 224806
<< end >>

