VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dcache
  CLASS BLOCK ;
  FOREIGN dcache ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 750.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END clk
  PIN d_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END d_in[0]
  PIN d_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END d_in[100]
  PIN d_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END d_in[101]
  PIN d_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END d_in[102]
  PIN d_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END d_in[103]
  PIN d_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END d_in[104]
  PIN d_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END d_in[105]
  PIN d_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END d_in[106]
  PIN d_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END d_in[107]
  PIN d_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END d_in[108]
  PIN d_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END d_in[109]
  PIN d_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END d_in[10]
  PIN d_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END d_in[110]
  PIN d_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END d_in[111]
  PIN d_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END d_in[112]
  PIN d_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END d_in[113]
  PIN d_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END d_in[114]
  PIN d_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END d_in[115]
  PIN d_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END d_in[116]
  PIN d_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END d_in[117]
  PIN d_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END d_in[118]
  PIN d_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END d_in[119]
  PIN d_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END d_in[11]
  PIN d_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END d_in[120]
  PIN d_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END d_in[121]
  PIN d_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END d_in[122]
  PIN d_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END d_in[123]
  PIN d_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END d_in[124]
  PIN d_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END d_in[125]
  PIN d_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END d_in[126]
  PIN d_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END d_in[127]
  PIN d_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END d_in[128]
  PIN d_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END d_in[129]
  PIN d_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END d_in[12]
  PIN d_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END d_in[130]
  PIN d_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END d_in[131]
  PIN d_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END d_in[132]
  PIN d_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END d_in[133]
  PIN d_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END d_in[134]
  PIN d_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END d_in[135]
  PIN d_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END d_in[136]
  PIN d_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END d_in[137]
  PIN d_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END d_in[138]
  PIN d_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END d_in[139]
  PIN d_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END d_in[13]
  PIN d_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END d_in[140]
  PIN d_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END d_in[141]
  PIN d_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END d_in[142]
  PIN d_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END d_in[14]
  PIN d_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END d_in[15]
  PIN d_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END d_in[16]
  PIN d_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END d_in[17]
  PIN d_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END d_in[18]
  PIN d_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END d_in[19]
  PIN d_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END d_in[1]
  PIN d_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END d_in[20]
  PIN d_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END d_in[21]
  PIN d_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END d_in[22]
  PIN d_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END d_in[23]
  PIN d_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END d_in[24]
  PIN d_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END d_in[25]
  PIN d_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END d_in[26]
  PIN d_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END d_in[27]
  PIN d_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END d_in[28]
  PIN d_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END d_in[29]
  PIN d_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END d_in[2]
  PIN d_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END d_in[30]
  PIN d_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END d_in[31]
  PIN d_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END d_in[32]
  PIN d_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END d_in[33]
  PIN d_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END d_in[34]
  PIN d_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END d_in[35]
  PIN d_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END d_in[36]
  PIN d_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END d_in[37]
  PIN d_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END d_in[38]
  PIN d_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END d_in[39]
  PIN d_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END d_in[3]
  PIN d_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END d_in[40]
  PIN d_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END d_in[41]
  PIN d_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END d_in[42]
  PIN d_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END d_in[43]
  PIN d_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END d_in[44]
  PIN d_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END d_in[45]
  PIN d_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END d_in[46]
  PIN d_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END d_in[47]
  PIN d_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END d_in[48]
  PIN d_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END d_in[49]
  PIN d_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END d_in[4]
  PIN d_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END d_in[50]
  PIN d_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END d_in[51]
  PIN d_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END d_in[52]
  PIN d_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END d_in[53]
  PIN d_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END d_in[54]
  PIN d_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END d_in[55]
  PIN d_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END d_in[56]
  PIN d_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END d_in[57]
  PIN d_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END d_in[58]
  PIN d_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END d_in[59]
  PIN d_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END d_in[5]
  PIN d_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END d_in[60]
  PIN d_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END d_in[61]
  PIN d_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END d_in[62]
  PIN d_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END d_in[63]
  PIN d_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END d_in[64]
  PIN d_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END d_in[65]
  PIN d_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END d_in[66]
  PIN d_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END d_in[67]
  PIN d_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END d_in[68]
  PIN d_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END d_in[69]
  PIN d_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END d_in[6]
  PIN d_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END d_in[70]
  PIN d_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END d_in[71]
  PIN d_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END d_in[72]
  PIN d_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END d_in[73]
  PIN d_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END d_in[74]
  PIN d_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END d_in[75]
  PIN d_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END d_in[76]
  PIN d_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END d_in[77]
  PIN d_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END d_in[78]
  PIN d_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END d_in[79]
  PIN d_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END d_in[7]
  PIN d_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END d_in[80]
  PIN d_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END d_in[81]
  PIN d_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END d_in[82]
  PIN d_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END d_in[83]
  PIN d_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END d_in[84]
  PIN d_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END d_in[85]
  PIN d_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END d_in[86]
  PIN d_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END d_in[87]
  PIN d_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END d_in[88]
  PIN d_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END d_in[89]
  PIN d_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END d_in[8]
  PIN d_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END d_in[90]
  PIN d_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END d_in[91]
  PIN d_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END d_in[92]
  PIN d_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END d_in[93]
  PIN d_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END d_in[94]
  PIN d_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END d_in[95]
  PIN d_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END d_in[96]
  PIN d_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END d_in[97]
  PIN d_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END d_in[98]
  PIN d_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END d_in[99]
  PIN d_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END d_in[9]
  PIN d_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END d_out[0]
  PIN d_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END d_out[10]
  PIN d_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END d_out[11]
  PIN d_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END d_out[12]
  PIN d_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END d_out[13]
  PIN d_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END d_out[14]
  PIN d_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END d_out[15]
  PIN d_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END d_out[16]
  PIN d_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END d_out[17]
  PIN d_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END d_out[18]
  PIN d_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END d_out[19]
  PIN d_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END d_out[1]
  PIN d_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END d_out[20]
  PIN d_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END d_out[21]
  PIN d_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END d_out[22]
  PIN d_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END d_out[23]
  PIN d_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END d_out[24]
  PIN d_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END d_out[25]
  PIN d_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END d_out[26]
  PIN d_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END d_out[27]
  PIN d_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END d_out[28]
  PIN d_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END d_out[29]
  PIN d_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END d_out[2]
  PIN d_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END d_out[30]
  PIN d_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END d_out[31]
  PIN d_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END d_out[32]
  PIN d_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 0.000 627.350 4.000 ;
    END
  END d_out[33]
  PIN d_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END d_out[34]
  PIN d_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END d_out[35]
  PIN d_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END d_out[36]
  PIN d_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END d_out[37]
  PIN d_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END d_out[38]
  PIN d_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END d_out[39]
  PIN d_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END d_out[3]
  PIN d_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END d_out[40]
  PIN d_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END d_out[41]
  PIN d_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 4.000 ;
    END
  END d_out[42]
  PIN d_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END d_out[43]
  PIN d_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END d_out[44]
  PIN d_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END d_out[45]
  PIN d_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END d_out[46]
  PIN d_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END d_out[47]
  PIN d_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END d_out[48]
  PIN d_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END d_out[49]
  PIN d_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END d_out[4]
  PIN d_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END d_out[50]
  PIN d_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END d_out[51]
  PIN d_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END d_out[52]
  PIN d_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END d_out[53]
  PIN d_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END d_out[54]
  PIN d_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END d_out[55]
  PIN d_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END d_out[56]
  PIN d_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END d_out[57]
  PIN d_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END d_out[58]
  PIN d_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END d_out[59]
  PIN d_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END d_out[5]
  PIN d_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END d_out[60]
  PIN d_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 4.000 ;
    END
  END d_out[61]
  PIN d_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END d_out[62]
  PIN d_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END d_out[63]
  PIN d_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END d_out[64]
  PIN d_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 0.000 740.510 4.000 ;
    END
  END d_out[65]
  PIN d_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END d_out[66]
  PIN d_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END d_out[67]
  PIN d_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END d_out[6]
  PIN d_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END d_out[7]
  PIN d_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END d_out[8]
  PIN d_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END d_out[9]
  PIN m_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END m_in[0]
  PIN m_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END m_in[100]
  PIN m_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END m_in[101]
  PIN m_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END m_in[102]
  PIN m_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END m_in[103]
  PIN m_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END m_in[104]
  PIN m_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.560 4.000 401.160 ;
    END
  END m_in[105]
  PIN m_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END m_in[106]
  PIN m_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END m_in[107]
  PIN m_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END m_in[108]
  PIN m_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END m_in[109]
  PIN m_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END m_in[10]
  PIN m_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END m_in[110]
  PIN m_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END m_in[111]
  PIN m_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END m_in[112]
  PIN m_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END m_in[113]
  PIN m_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END m_in[114]
  PIN m_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END m_in[115]
  PIN m_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END m_in[116]
  PIN m_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END m_in[117]
  PIN m_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END m_in[118]
  PIN m_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END m_in[119]
  PIN m_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END m_in[11]
  PIN m_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 4.000 456.920 ;
    END
  END m_in[120]
  PIN m_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END m_in[121]
  PIN m_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END m_in[122]
  PIN m_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.200 4.000 467.800 ;
    END
  END m_in[123]
  PIN m_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END m_in[124]
  PIN m_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END m_in[125]
  PIN m_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END m_in[126]
  PIN m_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END m_in[127]
  PIN m_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END m_in[128]
  PIN m_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END m_in[129]
  PIN m_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END m_in[12]
  PIN m_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END m_in[130]
  PIN m_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END m_in[131]
  PIN m_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END m_in[13]
  PIN m_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END m_in[14]
  PIN m_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END m_in[15]
  PIN m_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END m_in[16]
  PIN m_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END m_in[17]
  PIN m_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END m_in[18]
  PIN m_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END m_in[19]
  PIN m_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END m_in[1]
  PIN m_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END m_in[20]
  PIN m_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END m_in[21]
  PIN m_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END m_in[22]
  PIN m_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END m_in[23]
  PIN m_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END m_in[24]
  PIN m_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END m_in[25]
  PIN m_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END m_in[26]
  PIN m_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END m_in[27]
  PIN m_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END m_in[28]
  PIN m_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END m_in[29]
  PIN m_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END m_in[2]
  PIN m_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END m_in[30]
  PIN m_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END m_in[31]
  PIN m_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END m_in[32]
  PIN m_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END m_in[33]
  PIN m_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END m_in[34]
  PIN m_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END m_in[35]
  PIN m_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END m_in[36]
  PIN m_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END m_in[37]
  PIN m_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END m_in[38]
  PIN m_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END m_in[39]
  PIN m_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END m_in[3]
  PIN m_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END m_in[40]
  PIN m_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END m_in[41]
  PIN m_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END m_in[42]
  PIN m_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END m_in[43]
  PIN m_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END m_in[44]
  PIN m_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END m_in[45]
  PIN m_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END m_in[46]
  PIN m_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END m_in[47]
  PIN m_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END m_in[48]
  PIN m_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END m_in[49]
  PIN m_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END m_in[4]
  PIN m_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END m_in[50]
  PIN m_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END m_in[51]
  PIN m_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END m_in[52]
  PIN m_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END m_in[53]
  PIN m_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END m_in[54]
  PIN m_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END m_in[55]
  PIN m_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END m_in[56]
  PIN m_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END m_in[57]
  PIN m_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END m_in[58]
  PIN m_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END m_in[59]
  PIN m_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END m_in[5]
  PIN m_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END m_in[60]
  PIN m_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END m_in[61]
  PIN m_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END m_in[62]
  PIN m_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END m_in[63]
  PIN m_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END m_in[64]
  PIN m_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END m_in[65]
  PIN m_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END m_in[66]
  PIN m_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END m_in[67]
  PIN m_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END m_in[68]
  PIN m_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END m_in[69]
  PIN m_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END m_in[6]
  PIN m_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END m_in[70]
  PIN m_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END m_in[71]
  PIN m_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END m_in[72]
  PIN m_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END m_in[73]
  PIN m_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END m_in[74]
  PIN m_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END m_in[75]
  PIN m_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END m_in[76]
  PIN m_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END m_in[77]
  PIN m_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END m_in[78]
  PIN m_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END m_in[79]
  PIN m_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END m_in[7]
  PIN m_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END m_in[80]
  PIN m_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END m_in[81]
  PIN m_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END m_in[82]
  PIN m_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END m_in[83]
  PIN m_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END m_in[84]
  PIN m_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END m_in[85]
  PIN m_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END m_in[86]
  PIN m_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END m_in[87]
  PIN m_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END m_in[88]
  PIN m_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END m_in[89]
  PIN m_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END m_in[8]
  PIN m_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END m_in[90]
  PIN m_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END m_in[91]
  PIN m_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END m_in[92]
  PIN m_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END m_in[93]
  PIN m_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END m_in[94]
  PIN m_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END m_in[95]
  PIN m_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END m_in[96]
  PIN m_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END m_in[97]
  PIN m_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END m_in[98]
  PIN m_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END m_in[99]
  PIN m_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END m_in[9]
  PIN m_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END m_out[0]
  PIN m_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END m_out[10]
  PIN m_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END m_out[11]
  PIN m_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END m_out[12]
  PIN m_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END m_out[13]
  PIN m_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END m_out[14]
  PIN m_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END m_out[15]
  PIN m_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END m_out[16]
  PIN m_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END m_out[17]
  PIN m_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END m_out[18]
  PIN m_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END m_out[19]
  PIN m_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END m_out[1]
  PIN m_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.000 4.000 576.600 ;
    END
  END m_out[20]
  PIN m_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END m_out[21]
  PIN m_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END m_out[22]
  PIN m_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.880 4.000 587.480 ;
    END
  END m_out[23]
  PIN m_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END m_out[24]
  PIN m_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END m_out[25]
  PIN m_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END m_out[26]
  PIN m_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END m_out[27]
  PIN m_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END m_out[28]
  PIN m_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END m_out[29]
  PIN m_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END m_out[2]
  PIN m_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END m_out[30]
  PIN m_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END m_out[31]
  PIN m_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END m_out[32]
  PIN m_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END m_out[33]
  PIN m_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END m_out[34]
  PIN m_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END m_out[35]
  PIN m_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END m_out[36]
  PIN m_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END m_out[37]
  PIN m_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END m_out[38]
  PIN m_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END m_out[39]
  PIN m_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.080 4.000 512.680 ;
    END
  END m_out[3]
  PIN m_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END m_out[40]
  PIN m_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END m_out[41]
  PIN m_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END m_out[42]
  PIN m_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.680 4.000 662.280 ;
    END
  END m_out[43]
  PIN m_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END m_out[44]
  PIN m_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END m_out[45]
  PIN m_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 672.560 4.000 673.160 ;
    END
  END m_out[46]
  PIN m_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END m_out[47]
  PIN m_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END m_out[48]
  PIN m_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END m_out[49]
  PIN m_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.160 4.000 516.760 ;
    END
  END m_out[4]
  PIN m_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.520 4.000 688.120 ;
    END
  END m_out[50]
  PIN m_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END m_out[51]
  PIN m_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END m_out[52]
  PIN m_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END m_out[53]
  PIN m_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 702.480 4.000 703.080 ;
    END
  END m_out[54]
  PIN m_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 706.560 4.000 707.160 ;
    END
  END m_out[55]
  PIN m_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END m_out[56]
  PIN m_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END m_out[57]
  PIN m_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END m_out[58]
  PIN m_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 721.520 4.000 722.120 ;
    END
  END m_out[59]
  PIN m_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END m_out[5]
  PIN m_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END m_out[60]
  PIN m_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.000 4.000 729.600 ;
    END
  END m_out[61]
  PIN m_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 732.400 4.000 733.000 ;
    END
  END m_out[62]
  PIN m_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 736.480 4.000 737.080 ;
    END
  END m_out[63]
  PIN m_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END m_out[64]
  PIN m_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END m_out[65]
  PIN m_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 747.360 4.000 747.960 ;
    END
  END m_out[66]
  PIN m_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END m_out[6]
  PIN m_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END m_out[7]
  PIN m_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END m_out[8]
  PIN m_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END m_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END rst
  PIN stall_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END stall_out
  PIN wishbone_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 746.000 2.210 750.000 ;
    END
  END wishbone_in[0]
  PIN wishbone_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 746.000 45.450 750.000 ;
    END
  END wishbone_in[10]
  PIN wishbone_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 746.000 49.590 750.000 ;
    END
  END wishbone_in[11]
  PIN wishbone_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 746.000 54.190 750.000 ;
    END
  END wishbone_in[12]
  PIN wishbone_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 746.000 58.330 750.000 ;
    END
  END wishbone_in[13]
  PIN wishbone_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 746.000 62.470 750.000 ;
    END
  END wishbone_in[14]
  PIN wishbone_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 746.000 67.070 750.000 ;
    END
  END wishbone_in[15]
  PIN wishbone_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 746.000 71.210 750.000 ;
    END
  END wishbone_in[16]
  PIN wishbone_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 746.000 75.810 750.000 ;
    END
  END wishbone_in[17]
  PIN wishbone_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 746.000 79.950 750.000 ;
    END
  END wishbone_in[18]
  PIN wishbone_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 746.000 84.550 750.000 ;
    END
  END wishbone_in[19]
  PIN wishbone_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 746.000 6.350 750.000 ;
    END
  END wishbone_in[1]
  PIN wishbone_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 746.000 88.690 750.000 ;
    END
  END wishbone_in[20]
  PIN wishbone_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 746.000 92.830 750.000 ;
    END
  END wishbone_in[21]
  PIN wishbone_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 746.000 97.430 750.000 ;
    END
  END wishbone_in[22]
  PIN wishbone_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 746.000 101.570 750.000 ;
    END
  END wishbone_in[23]
  PIN wishbone_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 746.000 106.170 750.000 ;
    END
  END wishbone_in[24]
  PIN wishbone_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 746.000 110.310 750.000 ;
    END
  END wishbone_in[25]
  PIN wishbone_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 746.000 114.450 750.000 ;
    END
  END wishbone_in[26]
  PIN wishbone_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 746.000 119.050 750.000 ;
    END
  END wishbone_in[27]
  PIN wishbone_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 746.000 123.190 750.000 ;
    END
  END wishbone_in[28]
  PIN wishbone_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 746.000 127.790 750.000 ;
    END
  END wishbone_in[29]
  PIN wishbone_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 746.000 10.490 750.000 ;
    END
  END wishbone_in[2]
  PIN wishbone_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 746.000 131.930 750.000 ;
    END
  END wishbone_in[30]
  PIN wishbone_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 746.000 136.530 750.000 ;
    END
  END wishbone_in[31]
  PIN wishbone_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 746.000 140.670 750.000 ;
    END
  END wishbone_in[32]
  PIN wishbone_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 746.000 144.810 750.000 ;
    END
  END wishbone_in[33]
  PIN wishbone_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 746.000 149.410 750.000 ;
    END
  END wishbone_in[34]
  PIN wishbone_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 746.000 153.550 750.000 ;
    END
  END wishbone_in[35]
  PIN wishbone_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 746.000 158.150 750.000 ;
    END
  END wishbone_in[36]
  PIN wishbone_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 746.000 162.290 750.000 ;
    END
  END wishbone_in[37]
  PIN wishbone_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 746.000 166.890 750.000 ;
    END
  END wishbone_in[38]
  PIN wishbone_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 746.000 171.030 750.000 ;
    END
  END wishbone_in[39]
  PIN wishbone_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 746.000 15.090 750.000 ;
    END
  END wishbone_in[3]
  PIN wishbone_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 746.000 175.170 750.000 ;
    END
  END wishbone_in[40]
  PIN wishbone_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 746.000 179.770 750.000 ;
    END
  END wishbone_in[41]
  PIN wishbone_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 746.000 183.910 750.000 ;
    END
  END wishbone_in[42]
  PIN wishbone_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 746.000 188.510 750.000 ;
    END
  END wishbone_in[43]
  PIN wishbone_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 746.000 192.650 750.000 ;
    END
  END wishbone_in[44]
  PIN wishbone_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 746.000 196.790 750.000 ;
    END
  END wishbone_in[45]
  PIN wishbone_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 746.000 201.390 750.000 ;
    END
  END wishbone_in[46]
  PIN wishbone_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 746.000 205.530 750.000 ;
    END
  END wishbone_in[47]
  PIN wishbone_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 746.000 210.130 750.000 ;
    END
  END wishbone_in[48]
  PIN wishbone_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 746.000 214.270 750.000 ;
    END
  END wishbone_in[49]
  PIN wishbone_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 746.000 19.230 750.000 ;
    END
  END wishbone_in[4]
  PIN wishbone_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 746.000 218.870 750.000 ;
    END
  END wishbone_in[50]
  PIN wishbone_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 746.000 223.010 750.000 ;
    END
  END wishbone_in[51]
  PIN wishbone_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 746.000 227.150 750.000 ;
    END
  END wishbone_in[52]
  PIN wishbone_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 746.000 231.750 750.000 ;
    END
  END wishbone_in[53]
  PIN wishbone_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 746.000 235.890 750.000 ;
    END
  END wishbone_in[54]
  PIN wishbone_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 746.000 240.490 750.000 ;
    END
  END wishbone_in[55]
  PIN wishbone_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 746.000 244.630 750.000 ;
    END
  END wishbone_in[56]
  PIN wishbone_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 746.000 249.230 750.000 ;
    END
  END wishbone_in[57]
  PIN wishbone_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 746.000 253.370 750.000 ;
    END
  END wishbone_in[58]
  PIN wishbone_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 746.000 257.510 750.000 ;
    END
  END wishbone_in[59]
  PIN wishbone_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 746.000 23.830 750.000 ;
    END
  END wishbone_in[5]
  PIN wishbone_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 746.000 262.110 750.000 ;
    END
  END wishbone_in[60]
  PIN wishbone_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 746.000 266.250 750.000 ;
    END
  END wishbone_in[61]
  PIN wishbone_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 746.000 270.850 750.000 ;
    END
  END wishbone_in[62]
  PIN wishbone_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 746.000 274.990 750.000 ;
    END
  END wishbone_in[63]
  PIN wishbone_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 746.000 279.590 750.000 ;
    END
  END wishbone_in[64]
  PIN wishbone_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 746.000 283.730 750.000 ;
    END
  END wishbone_in[65]
  PIN wishbone_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 746.000 27.970 750.000 ;
    END
  END wishbone_in[6]
  PIN wishbone_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 746.000 32.110 750.000 ;
    END
  END wishbone_in[7]
  PIN wishbone_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 746.000 36.710 750.000 ;
    END
  END wishbone_in[8]
  PIN wishbone_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 746.000 40.850 750.000 ;
    END
  END wishbone_in[9]
  PIN wishbone_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 746.000 287.870 750.000 ;
    END
  END wishbone_out[0]
  PIN wishbone_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 746.000 721.650 750.000 ;
    END
  END wishbone_out[100]
  PIN wishbone_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 746.000 725.790 750.000 ;
    END
  END wishbone_out[101]
  PIN wishbone_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 746.000 729.930 750.000 ;
    END
  END wishbone_out[102]
  PIN wishbone_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 746.000 734.530 750.000 ;
    END
  END wishbone_out[103]
  PIN wishbone_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 746.000 738.670 750.000 ;
    END
  END wishbone_out[104]
  PIN wishbone_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 746.000 743.270 750.000 ;
    END
  END wishbone_out[105]
  PIN wishbone_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 746.000 747.410 750.000 ;
    END
  END wishbone_out[106]
  PIN wishbone_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 746.000 331.570 750.000 ;
    END
  END wishbone_out[10]
  PIN wishbone_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 746.000 335.710 750.000 ;
    END
  END wishbone_out[11]
  PIN wishbone_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 746.000 339.850 750.000 ;
    END
  END wishbone_out[12]
  PIN wishbone_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 746.000 344.450 750.000 ;
    END
  END wishbone_out[13]
  PIN wishbone_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 746.000 348.590 750.000 ;
    END
  END wishbone_out[14]
  PIN wishbone_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 746.000 353.190 750.000 ;
    END
  END wishbone_out[15]
  PIN wishbone_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 746.000 357.330 750.000 ;
    END
  END wishbone_out[16]
  PIN wishbone_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 746.000 361.930 750.000 ;
    END
  END wishbone_out[17]
  PIN wishbone_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 746.000 366.070 750.000 ;
    END
  END wishbone_out[18]
  PIN wishbone_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 746.000 370.210 750.000 ;
    END
  END wishbone_out[19]
  PIN wishbone_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 746.000 292.470 750.000 ;
    END
  END wishbone_out[1]
  PIN wishbone_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 746.000 374.810 750.000 ;
    END
  END wishbone_out[20]
  PIN wishbone_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 746.000 378.950 750.000 ;
    END
  END wishbone_out[21]
  PIN wishbone_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 746.000 383.550 750.000 ;
    END
  END wishbone_out[22]
  PIN wishbone_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 746.000 387.690 750.000 ;
    END
  END wishbone_out[23]
  PIN wishbone_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 746.000 391.830 750.000 ;
    END
  END wishbone_out[24]
  PIN wishbone_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 746.000 396.430 750.000 ;
    END
  END wishbone_out[25]
  PIN wishbone_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 746.000 400.570 750.000 ;
    END
  END wishbone_out[26]
  PIN wishbone_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 746.000 405.170 750.000 ;
    END
  END wishbone_out[27]
  PIN wishbone_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 746.000 409.310 750.000 ;
    END
  END wishbone_out[28]
  PIN wishbone_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 746.000 413.910 750.000 ;
    END
  END wishbone_out[29]
  PIN wishbone_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 746.000 296.610 750.000 ;
    END
  END wishbone_out[2]
  PIN wishbone_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 746.000 418.050 750.000 ;
    END
  END wishbone_out[30]
  PIN wishbone_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 746.000 422.190 750.000 ;
    END
  END wishbone_out[31]
  PIN wishbone_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 746.000 426.790 750.000 ;
    END
  END wishbone_out[32]
  PIN wishbone_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 746.000 430.930 750.000 ;
    END
  END wishbone_out[33]
  PIN wishbone_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 746.000 435.530 750.000 ;
    END
  END wishbone_out[34]
  PIN wishbone_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 746.000 439.670 750.000 ;
    END
  END wishbone_out[35]
  PIN wishbone_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 746.000 444.270 750.000 ;
    END
  END wishbone_out[36]
  PIN wishbone_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 746.000 448.410 750.000 ;
    END
  END wishbone_out[37]
  PIN wishbone_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 746.000 452.550 750.000 ;
    END
  END wishbone_out[38]
  PIN wishbone_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 746.000 457.150 750.000 ;
    END
  END wishbone_out[39]
  PIN wishbone_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 746.000 301.210 750.000 ;
    END
  END wishbone_out[3]
  PIN wishbone_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 746.000 461.290 750.000 ;
    END
  END wishbone_out[40]
  PIN wishbone_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 746.000 465.890 750.000 ;
    END
  END wishbone_out[41]
  PIN wishbone_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 746.000 470.030 750.000 ;
    END
  END wishbone_out[42]
  PIN wishbone_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 746.000 474.170 750.000 ;
    END
  END wishbone_out[43]
  PIN wishbone_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 746.000 478.770 750.000 ;
    END
  END wishbone_out[44]
  PIN wishbone_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 746.000 482.910 750.000 ;
    END
  END wishbone_out[45]
  PIN wishbone_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 746.000 487.510 750.000 ;
    END
  END wishbone_out[46]
  PIN wishbone_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 746.000 491.650 750.000 ;
    END
  END wishbone_out[47]
  PIN wishbone_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 746.000 496.250 750.000 ;
    END
  END wishbone_out[48]
  PIN wishbone_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 746.000 500.390 750.000 ;
    END
  END wishbone_out[49]
  PIN wishbone_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 746.000 305.350 750.000 ;
    END
  END wishbone_out[4]
  PIN wishbone_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 746.000 504.530 750.000 ;
    END
  END wishbone_out[50]
  PIN wishbone_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 746.000 509.130 750.000 ;
    END
  END wishbone_out[51]
  PIN wishbone_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 746.000 513.270 750.000 ;
    END
  END wishbone_out[52]
  PIN wishbone_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 746.000 517.870 750.000 ;
    END
  END wishbone_out[53]
  PIN wishbone_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 746.000 522.010 750.000 ;
    END
  END wishbone_out[54]
  PIN wishbone_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 746.000 526.610 750.000 ;
    END
  END wishbone_out[55]
  PIN wishbone_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 746.000 530.750 750.000 ;
    END
  END wishbone_out[56]
  PIN wishbone_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 746.000 534.890 750.000 ;
    END
  END wishbone_out[57]
  PIN wishbone_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 746.000 539.490 750.000 ;
    END
  END wishbone_out[58]
  PIN wishbone_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 746.000 543.630 750.000 ;
    END
  END wishbone_out[59]
  PIN wishbone_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 746.000 309.490 750.000 ;
    END
  END wishbone_out[5]
  PIN wishbone_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 746.000 548.230 750.000 ;
    END
  END wishbone_out[60]
  PIN wishbone_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 746.000 552.370 750.000 ;
    END
  END wishbone_out[61]
  PIN wishbone_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 746.000 556.970 750.000 ;
    END
  END wishbone_out[62]
  PIN wishbone_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 746.000 561.110 750.000 ;
    END
  END wishbone_out[63]
  PIN wishbone_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 746.000 565.250 750.000 ;
    END
  END wishbone_out[64]
  PIN wishbone_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 746.000 569.850 750.000 ;
    END
  END wishbone_out[65]
  PIN wishbone_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 746.000 573.990 750.000 ;
    END
  END wishbone_out[66]
  PIN wishbone_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 746.000 578.590 750.000 ;
    END
  END wishbone_out[67]
  PIN wishbone_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 746.000 582.730 750.000 ;
    END
  END wishbone_out[68]
  PIN wishbone_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 746.000 586.870 750.000 ;
    END
  END wishbone_out[69]
  PIN wishbone_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 746.000 314.090 750.000 ;
    END
  END wishbone_out[6]
  PIN wishbone_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 746.000 591.470 750.000 ;
    END
  END wishbone_out[70]
  PIN wishbone_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 746.000 595.610 750.000 ;
    END
  END wishbone_out[71]
  PIN wishbone_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 746.000 600.210 750.000 ;
    END
  END wishbone_out[72]
  PIN wishbone_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 746.000 604.350 750.000 ;
    END
  END wishbone_out[73]
  PIN wishbone_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 746.000 608.950 750.000 ;
    END
  END wishbone_out[74]
  PIN wishbone_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 746.000 613.090 750.000 ;
    END
  END wishbone_out[75]
  PIN wishbone_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 746.000 617.230 750.000 ;
    END
  END wishbone_out[76]
  PIN wishbone_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 746.000 621.830 750.000 ;
    END
  END wishbone_out[77]
  PIN wishbone_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 746.000 625.970 750.000 ;
    END
  END wishbone_out[78]
  PIN wishbone_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 746.000 630.570 750.000 ;
    END
  END wishbone_out[79]
  PIN wishbone_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 746.000 318.230 750.000 ;
    END
  END wishbone_out[7]
  PIN wishbone_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 746.000 634.710 750.000 ;
    END
  END wishbone_out[80]
  PIN wishbone_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 746.000 639.310 750.000 ;
    END
  END wishbone_out[81]
  PIN wishbone_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 746.000 643.450 750.000 ;
    END
  END wishbone_out[82]
  PIN wishbone_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 746.000 647.590 750.000 ;
    END
  END wishbone_out[83]
  PIN wishbone_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 746.000 652.190 750.000 ;
    END
  END wishbone_out[84]
  PIN wishbone_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 746.000 656.330 750.000 ;
    END
  END wishbone_out[85]
  PIN wishbone_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 746.000 660.930 750.000 ;
    END
  END wishbone_out[86]
  PIN wishbone_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 746.000 665.070 750.000 ;
    END
  END wishbone_out[87]
  PIN wishbone_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 746.000 669.210 750.000 ;
    END
  END wishbone_out[88]
  PIN wishbone_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 746.000 673.810 750.000 ;
    END
  END wishbone_out[89]
  PIN wishbone_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 746.000 322.830 750.000 ;
    END
  END wishbone_out[8]
  PIN wishbone_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 746.000 677.950 750.000 ;
    END
  END wishbone_out[90]
  PIN wishbone_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 746.000 682.550 750.000 ;
    END
  END wishbone_out[91]
  PIN wishbone_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 746.000 686.690 750.000 ;
    END
  END wishbone_out[92]
  PIN wishbone_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 746.000 691.290 750.000 ;
    END
  END wishbone_out[93]
  PIN wishbone_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 746.000 695.430 750.000 ;
    END
  END wishbone_out[94]
  PIN wishbone_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 746.000 699.570 750.000 ;
    END
  END wishbone_out[95]
  PIN wishbone_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 746.000 704.170 750.000 ;
    END
  END wishbone_out[96]
  PIN wishbone_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 746.000 708.310 750.000 ;
    END
  END wishbone_out[97]
  PIN wishbone_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 746.000 712.910 750.000 ;
    END
  END wishbone_out[98]
  PIN wishbone_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 746.000 717.050 750.000 ;
    END
  END wishbone_out[99]
  PIN wishbone_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 746.000 326.970 750.000 ;
    END
  END wishbone_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 737.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 737.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 737.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 737.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 737.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 737.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 737.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 737.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 737.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 737.360 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 744.280 737.205 ;
      LAYER met1 ;
        RECT 1.450 6.500 747.890 745.920 ;
      LAYER met2 ;
        RECT 1.480 745.720 1.650 747.845 ;
        RECT 2.490 745.720 5.790 747.845 ;
        RECT 6.630 745.720 9.930 747.845 ;
        RECT 10.770 745.720 14.530 747.845 ;
        RECT 15.370 745.720 18.670 747.845 ;
        RECT 19.510 745.720 23.270 747.845 ;
        RECT 24.110 745.720 27.410 747.845 ;
        RECT 28.250 745.720 31.550 747.845 ;
        RECT 32.390 745.720 36.150 747.845 ;
        RECT 36.990 745.720 40.290 747.845 ;
        RECT 41.130 745.720 44.890 747.845 ;
        RECT 45.730 745.720 49.030 747.845 ;
        RECT 49.870 745.720 53.630 747.845 ;
        RECT 54.470 745.720 57.770 747.845 ;
        RECT 58.610 745.720 61.910 747.845 ;
        RECT 62.750 745.720 66.510 747.845 ;
        RECT 67.350 745.720 70.650 747.845 ;
        RECT 71.490 745.720 75.250 747.845 ;
        RECT 76.090 745.720 79.390 747.845 ;
        RECT 80.230 745.720 83.990 747.845 ;
        RECT 84.830 745.720 88.130 747.845 ;
        RECT 88.970 745.720 92.270 747.845 ;
        RECT 93.110 745.720 96.870 747.845 ;
        RECT 97.710 745.720 101.010 747.845 ;
        RECT 101.850 745.720 105.610 747.845 ;
        RECT 106.450 745.720 109.750 747.845 ;
        RECT 110.590 745.720 113.890 747.845 ;
        RECT 114.730 745.720 118.490 747.845 ;
        RECT 119.330 745.720 122.630 747.845 ;
        RECT 123.470 745.720 127.230 747.845 ;
        RECT 128.070 745.720 131.370 747.845 ;
        RECT 132.210 745.720 135.970 747.845 ;
        RECT 136.810 745.720 140.110 747.845 ;
        RECT 140.950 745.720 144.250 747.845 ;
        RECT 145.090 745.720 148.850 747.845 ;
        RECT 149.690 745.720 152.990 747.845 ;
        RECT 153.830 745.720 157.590 747.845 ;
        RECT 158.430 745.720 161.730 747.845 ;
        RECT 162.570 745.720 166.330 747.845 ;
        RECT 167.170 745.720 170.470 747.845 ;
        RECT 171.310 745.720 174.610 747.845 ;
        RECT 175.450 745.720 179.210 747.845 ;
        RECT 180.050 745.720 183.350 747.845 ;
        RECT 184.190 745.720 187.950 747.845 ;
        RECT 188.790 745.720 192.090 747.845 ;
        RECT 192.930 745.720 196.230 747.845 ;
        RECT 197.070 745.720 200.830 747.845 ;
        RECT 201.670 745.720 204.970 747.845 ;
        RECT 205.810 745.720 209.570 747.845 ;
        RECT 210.410 745.720 213.710 747.845 ;
        RECT 214.550 745.720 218.310 747.845 ;
        RECT 219.150 745.720 222.450 747.845 ;
        RECT 223.290 745.720 226.590 747.845 ;
        RECT 227.430 745.720 231.190 747.845 ;
        RECT 232.030 745.720 235.330 747.845 ;
        RECT 236.170 745.720 239.930 747.845 ;
        RECT 240.770 745.720 244.070 747.845 ;
        RECT 244.910 745.720 248.670 747.845 ;
        RECT 249.510 745.720 252.810 747.845 ;
        RECT 253.650 745.720 256.950 747.845 ;
        RECT 257.790 745.720 261.550 747.845 ;
        RECT 262.390 745.720 265.690 747.845 ;
        RECT 266.530 745.720 270.290 747.845 ;
        RECT 271.130 745.720 274.430 747.845 ;
        RECT 275.270 745.720 279.030 747.845 ;
        RECT 279.870 745.720 283.170 747.845 ;
        RECT 284.010 745.720 287.310 747.845 ;
        RECT 288.150 745.720 291.910 747.845 ;
        RECT 292.750 745.720 296.050 747.845 ;
        RECT 296.890 745.720 300.650 747.845 ;
        RECT 301.490 745.720 304.790 747.845 ;
        RECT 305.630 745.720 308.930 747.845 ;
        RECT 309.770 745.720 313.530 747.845 ;
        RECT 314.370 745.720 317.670 747.845 ;
        RECT 318.510 745.720 322.270 747.845 ;
        RECT 323.110 745.720 326.410 747.845 ;
        RECT 327.250 745.720 331.010 747.845 ;
        RECT 331.850 745.720 335.150 747.845 ;
        RECT 335.990 745.720 339.290 747.845 ;
        RECT 340.130 745.720 343.890 747.845 ;
        RECT 344.730 745.720 348.030 747.845 ;
        RECT 348.870 745.720 352.630 747.845 ;
        RECT 353.470 745.720 356.770 747.845 ;
        RECT 357.610 745.720 361.370 747.845 ;
        RECT 362.210 745.720 365.510 747.845 ;
        RECT 366.350 745.720 369.650 747.845 ;
        RECT 370.490 745.720 374.250 747.845 ;
        RECT 375.090 745.720 378.390 747.845 ;
        RECT 379.230 745.720 382.990 747.845 ;
        RECT 383.830 745.720 387.130 747.845 ;
        RECT 387.970 745.720 391.270 747.845 ;
        RECT 392.110 745.720 395.870 747.845 ;
        RECT 396.710 745.720 400.010 747.845 ;
        RECT 400.850 745.720 404.610 747.845 ;
        RECT 405.450 745.720 408.750 747.845 ;
        RECT 409.590 745.720 413.350 747.845 ;
        RECT 414.190 745.720 417.490 747.845 ;
        RECT 418.330 745.720 421.630 747.845 ;
        RECT 422.470 745.720 426.230 747.845 ;
        RECT 427.070 745.720 430.370 747.845 ;
        RECT 431.210 745.720 434.970 747.845 ;
        RECT 435.810 745.720 439.110 747.845 ;
        RECT 439.950 745.720 443.710 747.845 ;
        RECT 444.550 745.720 447.850 747.845 ;
        RECT 448.690 745.720 451.990 747.845 ;
        RECT 452.830 745.720 456.590 747.845 ;
        RECT 457.430 745.720 460.730 747.845 ;
        RECT 461.570 745.720 465.330 747.845 ;
        RECT 466.170 745.720 469.470 747.845 ;
        RECT 470.310 745.720 473.610 747.845 ;
        RECT 474.450 745.720 478.210 747.845 ;
        RECT 479.050 745.720 482.350 747.845 ;
        RECT 483.190 745.720 486.950 747.845 ;
        RECT 487.790 745.720 491.090 747.845 ;
        RECT 491.930 745.720 495.690 747.845 ;
        RECT 496.530 745.720 499.830 747.845 ;
        RECT 500.670 745.720 503.970 747.845 ;
        RECT 504.810 745.720 508.570 747.845 ;
        RECT 509.410 745.720 512.710 747.845 ;
        RECT 513.550 745.720 517.310 747.845 ;
        RECT 518.150 745.720 521.450 747.845 ;
        RECT 522.290 745.720 526.050 747.845 ;
        RECT 526.890 745.720 530.190 747.845 ;
        RECT 531.030 745.720 534.330 747.845 ;
        RECT 535.170 745.720 538.930 747.845 ;
        RECT 539.770 745.720 543.070 747.845 ;
        RECT 543.910 745.720 547.670 747.845 ;
        RECT 548.510 745.720 551.810 747.845 ;
        RECT 552.650 745.720 556.410 747.845 ;
        RECT 557.250 745.720 560.550 747.845 ;
        RECT 561.390 745.720 564.690 747.845 ;
        RECT 565.530 745.720 569.290 747.845 ;
        RECT 570.130 745.720 573.430 747.845 ;
        RECT 574.270 745.720 578.030 747.845 ;
        RECT 578.870 745.720 582.170 747.845 ;
        RECT 583.010 745.720 586.310 747.845 ;
        RECT 587.150 745.720 590.910 747.845 ;
        RECT 591.750 745.720 595.050 747.845 ;
        RECT 595.890 745.720 599.650 747.845 ;
        RECT 600.490 745.720 603.790 747.845 ;
        RECT 604.630 745.720 608.390 747.845 ;
        RECT 609.230 745.720 612.530 747.845 ;
        RECT 613.370 745.720 616.670 747.845 ;
        RECT 617.510 745.720 621.270 747.845 ;
        RECT 622.110 745.720 625.410 747.845 ;
        RECT 626.250 745.720 630.010 747.845 ;
        RECT 630.850 745.720 634.150 747.845 ;
        RECT 634.990 745.720 638.750 747.845 ;
        RECT 639.590 745.720 642.890 747.845 ;
        RECT 643.730 745.720 647.030 747.845 ;
        RECT 647.870 745.720 651.630 747.845 ;
        RECT 652.470 745.720 655.770 747.845 ;
        RECT 656.610 745.720 660.370 747.845 ;
        RECT 661.210 745.720 664.510 747.845 ;
        RECT 665.350 745.720 668.650 747.845 ;
        RECT 669.490 745.720 673.250 747.845 ;
        RECT 674.090 745.720 677.390 747.845 ;
        RECT 678.230 745.720 681.990 747.845 ;
        RECT 682.830 745.720 686.130 747.845 ;
        RECT 686.970 745.720 690.730 747.845 ;
        RECT 691.570 745.720 694.870 747.845 ;
        RECT 695.710 745.720 699.010 747.845 ;
        RECT 699.850 745.720 703.610 747.845 ;
        RECT 704.450 745.720 707.750 747.845 ;
        RECT 708.590 745.720 712.350 747.845 ;
        RECT 713.190 745.720 716.490 747.845 ;
        RECT 717.330 745.720 721.090 747.845 ;
        RECT 721.930 745.720 725.230 747.845 ;
        RECT 726.070 745.720 729.370 747.845 ;
        RECT 730.210 745.720 733.970 747.845 ;
        RECT 734.810 745.720 738.110 747.845 ;
        RECT 738.950 745.720 742.710 747.845 ;
        RECT 743.550 745.720 746.850 747.845 ;
        RECT 747.690 745.720 747.860 747.845 ;
        RECT 1.480 4.280 747.860 745.720 ;
        RECT 2.030 1.515 4.410 4.280 ;
        RECT 5.250 1.515 8.090 4.280 ;
        RECT 8.930 1.515 11.770 4.280 ;
        RECT 12.610 1.515 14.990 4.280 ;
        RECT 15.830 1.515 18.670 4.280 ;
        RECT 19.510 1.515 22.350 4.280 ;
        RECT 23.190 1.515 25.570 4.280 ;
        RECT 26.410 1.515 29.250 4.280 ;
        RECT 30.090 1.515 32.930 4.280 ;
        RECT 33.770 1.515 36.150 4.280 ;
        RECT 36.990 1.515 39.830 4.280 ;
        RECT 40.670 1.515 43.510 4.280 ;
        RECT 44.350 1.515 46.730 4.280 ;
        RECT 47.570 1.515 50.410 4.280 ;
        RECT 51.250 1.515 54.090 4.280 ;
        RECT 54.930 1.515 57.770 4.280 ;
        RECT 58.610 1.515 60.990 4.280 ;
        RECT 61.830 1.515 64.670 4.280 ;
        RECT 65.510 1.515 68.350 4.280 ;
        RECT 69.190 1.515 71.570 4.280 ;
        RECT 72.410 1.515 75.250 4.280 ;
        RECT 76.090 1.515 78.930 4.280 ;
        RECT 79.770 1.515 82.150 4.280 ;
        RECT 82.990 1.515 85.830 4.280 ;
        RECT 86.670 1.515 89.510 4.280 ;
        RECT 90.350 1.515 92.730 4.280 ;
        RECT 93.570 1.515 96.410 4.280 ;
        RECT 97.250 1.515 100.090 4.280 ;
        RECT 100.930 1.515 103.310 4.280 ;
        RECT 104.150 1.515 106.990 4.280 ;
        RECT 107.830 1.515 110.670 4.280 ;
        RECT 111.510 1.515 114.350 4.280 ;
        RECT 115.190 1.515 117.570 4.280 ;
        RECT 118.410 1.515 121.250 4.280 ;
        RECT 122.090 1.515 124.930 4.280 ;
        RECT 125.770 1.515 128.150 4.280 ;
        RECT 128.990 1.515 131.830 4.280 ;
        RECT 132.670 1.515 135.510 4.280 ;
        RECT 136.350 1.515 138.730 4.280 ;
        RECT 139.570 1.515 142.410 4.280 ;
        RECT 143.250 1.515 146.090 4.280 ;
        RECT 146.930 1.515 149.310 4.280 ;
        RECT 150.150 1.515 152.990 4.280 ;
        RECT 153.830 1.515 156.670 4.280 ;
        RECT 157.510 1.515 159.890 4.280 ;
        RECT 160.730 1.515 163.570 4.280 ;
        RECT 164.410 1.515 167.250 4.280 ;
        RECT 168.090 1.515 170.930 4.280 ;
        RECT 171.770 1.515 174.150 4.280 ;
        RECT 174.990 1.515 177.830 4.280 ;
        RECT 178.670 1.515 181.510 4.280 ;
        RECT 182.350 1.515 184.730 4.280 ;
        RECT 185.570 1.515 188.410 4.280 ;
        RECT 189.250 1.515 192.090 4.280 ;
        RECT 192.930 1.515 195.310 4.280 ;
        RECT 196.150 1.515 198.990 4.280 ;
        RECT 199.830 1.515 202.670 4.280 ;
        RECT 203.510 1.515 205.890 4.280 ;
        RECT 206.730 1.515 209.570 4.280 ;
        RECT 210.410 1.515 213.250 4.280 ;
        RECT 214.090 1.515 216.930 4.280 ;
        RECT 217.770 1.515 220.150 4.280 ;
        RECT 220.990 1.515 223.830 4.280 ;
        RECT 224.670 1.515 227.510 4.280 ;
        RECT 228.350 1.515 230.730 4.280 ;
        RECT 231.570 1.515 234.410 4.280 ;
        RECT 235.250 1.515 238.090 4.280 ;
        RECT 238.930 1.515 241.310 4.280 ;
        RECT 242.150 1.515 244.990 4.280 ;
        RECT 245.830 1.515 248.670 4.280 ;
        RECT 249.510 1.515 251.890 4.280 ;
        RECT 252.730 1.515 255.570 4.280 ;
        RECT 256.410 1.515 259.250 4.280 ;
        RECT 260.090 1.515 262.470 4.280 ;
        RECT 263.310 1.515 266.150 4.280 ;
        RECT 266.990 1.515 269.830 4.280 ;
        RECT 270.670 1.515 273.510 4.280 ;
        RECT 274.350 1.515 276.730 4.280 ;
        RECT 277.570 1.515 280.410 4.280 ;
        RECT 281.250 1.515 284.090 4.280 ;
        RECT 284.930 1.515 287.310 4.280 ;
        RECT 288.150 1.515 290.990 4.280 ;
        RECT 291.830 1.515 294.670 4.280 ;
        RECT 295.510 1.515 297.890 4.280 ;
        RECT 298.730 1.515 301.570 4.280 ;
        RECT 302.410 1.515 305.250 4.280 ;
        RECT 306.090 1.515 308.470 4.280 ;
        RECT 309.310 1.515 312.150 4.280 ;
        RECT 312.990 1.515 315.830 4.280 ;
        RECT 316.670 1.515 319.050 4.280 ;
        RECT 319.890 1.515 322.730 4.280 ;
        RECT 323.570 1.515 326.410 4.280 ;
        RECT 327.250 1.515 330.090 4.280 ;
        RECT 330.930 1.515 333.310 4.280 ;
        RECT 334.150 1.515 336.990 4.280 ;
        RECT 337.830 1.515 340.670 4.280 ;
        RECT 341.510 1.515 343.890 4.280 ;
        RECT 344.730 1.515 347.570 4.280 ;
        RECT 348.410 1.515 351.250 4.280 ;
        RECT 352.090 1.515 354.470 4.280 ;
        RECT 355.310 1.515 358.150 4.280 ;
        RECT 358.990 1.515 361.830 4.280 ;
        RECT 362.670 1.515 365.050 4.280 ;
        RECT 365.890 1.515 368.730 4.280 ;
        RECT 369.570 1.515 372.410 4.280 ;
        RECT 373.250 1.515 376.090 4.280 ;
        RECT 376.930 1.515 379.310 4.280 ;
        RECT 380.150 1.515 382.990 4.280 ;
        RECT 383.830 1.515 386.670 4.280 ;
        RECT 387.510 1.515 389.890 4.280 ;
        RECT 390.730 1.515 393.570 4.280 ;
        RECT 394.410 1.515 397.250 4.280 ;
        RECT 398.090 1.515 400.470 4.280 ;
        RECT 401.310 1.515 404.150 4.280 ;
        RECT 404.990 1.515 407.830 4.280 ;
        RECT 408.670 1.515 411.050 4.280 ;
        RECT 411.890 1.515 414.730 4.280 ;
        RECT 415.570 1.515 418.410 4.280 ;
        RECT 419.250 1.515 421.630 4.280 ;
        RECT 422.470 1.515 425.310 4.280 ;
        RECT 426.150 1.515 428.990 4.280 ;
        RECT 429.830 1.515 432.670 4.280 ;
        RECT 433.510 1.515 435.890 4.280 ;
        RECT 436.730 1.515 439.570 4.280 ;
        RECT 440.410 1.515 443.250 4.280 ;
        RECT 444.090 1.515 446.470 4.280 ;
        RECT 447.310 1.515 450.150 4.280 ;
        RECT 450.990 1.515 453.830 4.280 ;
        RECT 454.670 1.515 457.050 4.280 ;
        RECT 457.890 1.515 460.730 4.280 ;
        RECT 461.570 1.515 464.410 4.280 ;
        RECT 465.250 1.515 467.630 4.280 ;
        RECT 468.470 1.515 471.310 4.280 ;
        RECT 472.150 1.515 474.990 4.280 ;
        RECT 475.830 1.515 478.210 4.280 ;
        RECT 479.050 1.515 481.890 4.280 ;
        RECT 482.730 1.515 485.570 4.280 ;
        RECT 486.410 1.515 489.250 4.280 ;
        RECT 490.090 1.515 492.470 4.280 ;
        RECT 493.310 1.515 496.150 4.280 ;
        RECT 496.990 1.515 499.830 4.280 ;
        RECT 500.670 1.515 503.050 4.280 ;
        RECT 503.890 1.515 506.730 4.280 ;
        RECT 507.570 1.515 510.410 4.280 ;
        RECT 511.250 1.515 513.630 4.280 ;
        RECT 514.470 1.515 517.310 4.280 ;
        RECT 518.150 1.515 520.990 4.280 ;
        RECT 521.830 1.515 524.210 4.280 ;
        RECT 525.050 1.515 527.890 4.280 ;
        RECT 528.730 1.515 531.570 4.280 ;
        RECT 532.410 1.515 534.790 4.280 ;
        RECT 535.630 1.515 538.470 4.280 ;
        RECT 539.310 1.515 542.150 4.280 ;
        RECT 542.990 1.515 545.830 4.280 ;
        RECT 546.670 1.515 549.050 4.280 ;
        RECT 549.890 1.515 552.730 4.280 ;
        RECT 553.570 1.515 556.410 4.280 ;
        RECT 557.250 1.515 559.630 4.280 ;
        RECT 560.470 1.515 563.310 4.280 ;
        RECT 564.150 1.515 566.990 4.280 ;
        RECT 567.830 1.515 570.210 4.280 ;
        RECT 571.050 1.515 573.890 4.280 ;
        RECT 574.730 1.515 577.570 4.280 ;
        RECT 578.410 1.515 580.790 4.280 ;
        RECT 581.630 1.515 584.470 4.280 ;
        RECT 585.310 1.515 588.150 4.280 ;
        RECT 588.990 1.515 591.830 4.280 ;
        RECT 592.670 1.515 595.050 4.280 ;
        RECT 595.890 1.515 598.730 4.280 ;
        RECT 599.570 1.515 602.410 4.280 ;
        RECT 603.250 1.515 605.630 4.280 ;
        RECT 606.470 1.515 609.310 4.280 ;
        RECT 610.150 1.515 612.990 4.280 ;
        RECT 613.830 1.515 616.210 4.280 ;
        RECT 617.050 1.515 619.890 4.280 ;
        RECT 620.730 1.515 623.570 4.280 ;
        RECT 624.410 1.515 626.790 4.280 ;
        RECT 627.630 1.515 630.470 4.280 ;
        RECT 631.310 1.515 634.150 4.280 ;
        RECT 634.990 1.515 637.370 4.280 ;
        RECT 638.210 1.515 641.050 4.280 ;
        RECT 641.890 1.515 644.730 4.280 ;
        RECT 645.570 1.515 648.410 4.280 ;
        RECT 649.250 1.515 651.630 4.280 ;
        RECT 652.470 1.515 655.310 4.280 ;
        RECT 656.150 1.515 658.990 4.280 ;
        RECT 659.830 1.515 662.210 4.280 ;
        RECT 663.050 1.515 665.890 4.280 ;
        RECT 666.730 1.515 669.570 4.280 ;
        RECT 670.410 1.515 672.790 4.280 ;
        RECT 673.630 1.515 676.470 4.280 ;
        RECT 677.310 1.515 680.150 4.280 ;
        RECT 680.990 1.515 683.370 4.280 ;
        RECT 684.210 1.515 687.050 4.280 ;
        RECT 687.890 1.515 690.730 4.280 ;
        RECT 691.570 1.515 693.950 4.280 ;
        RECT 694.790 1.515 697.630 4.280 ;
        RECT 698.470 1.515 701.310 4.280 ;
        RECT 702.150 1.515 704.990 4.280 ;
        RECT 705.830 1.515 708.210 4.280 ;
        RECT 709.050 1.515 711.890 4.280 ;
        RECT 712.730 1.515 715.570 4.280 ;
        RECT 716.410 1.515 718.790 4.280 ;
        RECT 719.630 1.515 722.470 4.280 ;
        RECT 723.310 1.515 726.150 4.280 ;
        RECT 726.990 1.515 729.370 4.280 ;
        RECT 730.210 1.515 733.050 4.280 ;
        RECT 733.890 1.515 736.730 4.280 ;
        RECT 737.570 1.515 739.950 4.280 ;
        RECT 740.790 1.515 743.630 4.280 ;
        RECT 744.470 1.515 747.310 4.280 ;
      LAYER met3 ;
        RECT 4.400 746.960 741.915 747.825 ;
        RECT 1.190 744.960 741.915 746.960 ;
        RECT 4.400 743.560 741.915 744.960 ;
        RECT 1.190 740.880 741.915 743.560 ;
        RECT 4.400 739.480 741.915 740.880 ;
        RECT 1.190 737.480 741.915 739.480 ;
        RECT 4.400 736.080 741.915 737.480 ;
        RECT 1.190 733.400 741.915 736.080 ;
        RECT 4.400 732.000 741.915 733.400 ;
        RECT 1.190 730.000 741.915 732.000 ;
        RECT 4.400 728.600 741.915 730.000 ;
        RECT 1.190 725.920 741.915 728.600 ;
        RECT 4.400 724.520 741.915 725.920 ;
        RECT 1.190 722.520 741.915 724.520 ;
        RECT 4.400 721.120 741.915 722.520 ;
        RECT 1.190 718.440 741.915 721.120 ;
        RECT 4.400 717.040 741.915 718.440 ;
        RECT 1.190 715.040 741.915 717.040 ;
        RECT 4.400 713.640 741.915 715.040 ;
        RECT 1.190 710.960 741.915 713.640 ;
        RECT 4.400 709.560 741.915 710.960 ;
        RECT 1.190 707.560 741.915 709.560 ;
        RECT 4.400 706.160 741.915 707.560 ;
        RECT 1.190 703.480 741.915 706.160 ;
        RECT 4.400 702.080 741.915 703.480 ;
        RECT 1.190 700.080 741.915 702.080 ;
        RECT 4.400 698.680 741.915 700.080 ;
        RECT 1.190 696.000 741.915 698.680 ;
        RECT 4.400 694.600 741.915 696.000 ;
        RECT 1.190 692.600 741.915 694.600 ;
        RECT 4.400 691.200 741.915 692.600 ;
        RECT 1.190 688.520 741.915 691.200 ;
        RECT 4.400 687.120 741.915 688.520 ;
        RECT 1.190 685.120 741.915 687.120 ;
        RECT 4.400 683.720 741.915 685.120 ;
        RECT 1.190 681.040 741.915 683.720 ;
        RECT 4.400 679.640 741.915 681.040 ;
        RECT 1.190 677.640 741.915 679.640 ;
        RECT 4.400 676.240 741.915 677.640 ;
        RECT 1.190 673.560 741.915 676.240 ;
        RECT 4.400 672.160 741.915 673.560 ;
        RECT 1.190 670.160 741.915 672.160 ;
        RECT 4.400 668.760 741.915 670.160 ;
        RECT 1.190 666.080 741.915 668.760 ;
        RECT 4.400 664.680 741.915 666.080 ;
        RECT 1.190 662.680 741.915 664.680 ;
        RECT 4.400 661.280 741.915 662.680 ;
        RECT 1.190 658.600 741.915 661.280 ;
        RECT 4.400 657.200 741.915 658.600 ;
        RECT 1.190 655.200 741.915 657.200 ;
        RECT 4.400 653.800 741.915 655.200 ;
        RECT 1.190 651.120 741.915 653.800 ;
        RECT 4.400 649.720 741.915 651.120 ;
        RECT 1.190 647.720 741.915 649.720 ;
        RECT 4.400 646.320 741.915 647.720 ;
        RECT 1.190 643.640 741.915 646.320 ;
        RECT 4.400 642.240 741.915 643.640 ;
        RECT 1.190 640.240 741.915 642.240 ;
        RECT 4.400 638.840 741.915 640.240 ;
        RECT 1.190 636.160 741.915 638.840 ;
        RECT 4.400 634.760 741.915 636.160 ;
        RECT 1.190 632.760 741.915 634.760 ;
        RECT 4.400 631.360 741.915 632.760 ;
        RECT 1.190 628.680 741.915 631.360 ;
        RECT 4.400 627.280 741.915 628.680 ;
        RECT 1.190 625.280 741.915 627.280 ;
        RECT 4.400 623.880 741.915 625.280 ;
        RECT 1.190 621.200 741.915 623.880 ;
        RECT 4.400 619.800 741.915 621.200 ;
        RECT 1.190 617.800 741.915 619.800 ;
        RECT 4.400 616.400 741.915 617.800 ;
        RECT 1.190 613.720 741.915 616.400 ;
        RECT 4.400 612.320 741.915 613.720 ;
        RECT 1.190 610.320 741.915 612.320 ;
        RECT 4.400 608.920 741.915 610.320 ;
        RECT 1.190 606.240 741.915 608.920 ;
        RECT 4.400 604.840 741.915 606.240 ;
        RECT 1.190 602.840 741.915 604.840 ;
        RECT 4.400 601.440 741.915 602.840 ;
        RECT 1.190 599.440 741.915 601.440 ;
        RECT 4.400 598.040 741.915 599.440 ;
        RECT 1.190 595.360 741.915 598.040 ;
        RECT 4.400 593.960 741.915 595.360 ;
        RECT 1.190 591.960 741.915 593.960 ;
        RECT 4.400 590.560 741.915 591.960 ;
        RECT 1.190 587.880 741.915 590.560 ;
        RECT 4.400 586.480 741.915 587.880 ;
        RECT 1.190 584.480 741.915 586.480 ;
        RECT 4.400 583.080 741.915 584.480 ;
        RECT 1.190 580.400 741.915 583.080 ;
        RECT 4.400 579.000 741.915 580.400 ;
        RECT 1.190 577.000 741.915 579.000 ;
        RECT 4.400 575.600 741.915 577.000 ;
        RECT 1.190 572.920 741.915 575.600 ;
        RECT 4.400 571.520 741.915 572.920 ;
        RECT 1.190 569.520 741.915 571.520 ;
        RECT 4.400 568.120 741.915 569.520 ;
        RECT 1.190 565.440 741.915 568.120 ;
        RECT 4.400 564.040 741.915 565.440 ;
        RECT 1.190 562.040 741.915 564.040 ;
        RECT 4.400 560.640 741.915 562.040 ;
        RECT 1.190 557.960 741.915 560.640 ;
        RECT 4.400 556.560 741.915 557.960 ;
        RECT 1.190 554.560 741.915 556.560 ;
        RECT 4.400 553.160 741.915 554.560 ;
        RECT 1.190 550.480 741.915 553.160 ;
        RECT 4.400 549.080 741.915 550.480 ;
        RECT 1.190 547.080 741.915 549.080 ;
        RECT 4.400 545.680 741.915 547.080 ;
        RECT 1.190 543.000 741.915 545.680 ;
        RECT 4.400 541.600 741.915 543.000 ;
        RECT 1.190 539.600 741.915 541.600 ;
        RECT 4.400 538.200 741.915 539.600 ;
        RECT 1.190 535.520 741.915 538.200 ;
        RECT 4.400 534.120 741.915 535.520 ;
        RECT 1.190 532.120 741.915 534.120 ;
        RECT 4.400 530.720 741.915 532.120 ;
        RECT 1.190 528.040 741.915 530.720 ;
        RECT 4.400 526.640 741.915 528.040 ;
        RECT 1.190 524.640 741.915 526.640 ;
        RECT 4.400 523.240 741.915 524.640 ;
        RECT 1.190 520.560 741.915 523.240 ;
        RECT 4.400 519.160 741.915 520.560 ;
        RECT 1.190 517.160 741.915 519.160 ;
        RECT 4.400 515.760 741.915 517.160 ;
        RECT 1.190 513.080 741.915 515.760 ;
        RECT 4.400 511.680 741.915 513.080 ;
        RECT 1.190 509.680 741.915 511.680 ;
        RECT 4.400 508.280 741.915 509.680 ;
        RECT 1.190 505.600 741.915 508.280 ;
        RECT 4.400 504.200 741.915 505.600 ;
        RECT 1.190 502.200 741.915 504.200 ;
        RECT 4.400 500.800 741.915 502.200 ;
        RECT 1.190 498.120 741.915 500.800 ;
        RECT 4.400 496.720 741.915 498.120 ;
        RECT 1.190 494.720 741.915 496.720 ;
        RECT 4.400 493.320 741.915 494.720 ;
        RECT 1.190 490.640 741.915 493.320 ;
        RECT 4.400 489.240 741.915 490.640 ;
        RECT 1.190 487.240 741.915 489.240 ;
        RECT 4.400 485.840 741.915 487.240 ;
        RECT 1.190 483.160 741.915 485.840 ;
        RECT 4.400 481.760 741.915 483.160 ;
        RECT 1.190 479.760 741.915 481.760 ;
        RECT 4.400 478.360 741.915 479.760 ;
        RECT 1.190 475.680 741.915 478.360 ;
        RECT 4.400 474.280 741.915 475.680 ;
        RECT 1.190 472.280 741.915 474.280 ;
        RECT 4.400 470.880 741.915 472.280 ;
        RECT 1.190 468.200 741.915 470.880 ;
        RECT 4.400 466.800 741.915 468.200 ;
        RECT 1.190 464.800 741.915 466.800 ;
        RECT 4.400 463.400 741.915 464.800 ;
        RECT 1.190 460.720 741.915 463.400 ;
        RECT 4.400 459.320 741.915 460.720 ;
        RECT 1.190 457.320 741.915 459.320 ;
        RECT 4.400 455.920 741.915 457.320 ;
        RECT 1.190 453.240 741.915 455.920 ;
        RECT 4.400 451.840 741.915 453.240 ;
        RECT 1.190 449.840 741.915 451.840 ;
        RECT 4.400 448.440 741.915 449.840 ;
        RECT 1.190 446.440 741.915 448.440 ;
        RECT 4.400 445.040 741.915 446.440 ;
        RECT 1.190 442.360 741.915 445.040 ;
        RECT 4.400 440.960 741.915 442.360 ;
        RECT 1.190 438.960 741.915 440.960 ;
        RECT 4.400 437.560 741.915 438.960 ;
        RECT 1.190 434.880 741.915 437.560 ;
        RECT 4.400 433.480 741.915 434.880 ;
        RECT 1.190 431.480 741.915 433.480 ;
        RECT 4.400 430.080 741.915 431.480 ;
        RECT 1.190 427.400 741.915 430.080 ;
        RECT 4.400 426.000 741.915 427.400 ;
        RECT 1.190 424.000 741.915 426.000 ;
        RECT 4.400 422.600 741.915 424.000 ;
        RECT 1.190 419.920 741.915 422.600 ;
        RECT 4.400 418.520 741.915 419.920 ;
        RECT 1.190 416.520 741.915 418.520 ;
        RECT 4.400 415.120 741.915 416.520 ;
        RECT 1.190 412.440 741.915 415.120 ;
        RECT 4.400 411.040 741.915 412.440 ;
        RECT 1.190 409.040 741.915 411.040 ;
        RECT 4.400 407.640 741.915 409.040 ;
        RECT 1.190 404.960 741.915 407.640 ;
        RECT 4.400 403.560 741.915 404.960 ;
        RECT 1.190 401.560 741.915 403.560 ;
        RECT 4.400 400.160 741.915 401.560 ;
        RECT 1.190 397.480 741.915 400.160 ;
        RECT 4.400 396.080 741.915 397.480 ;
        RECT 1.190 394.080 741.915 396.080 ;
        RECT 4.400 392.680 741.915 394.080 ;
        RECT 1.190 390.000 741.915 392.680 ;
        RECT 4.400 388.600 741.915 390.000 ;
        RECT 1.190 386.600 741.915 388.600 ;
        RECT 4.400 385.200 741.915 386.600 ;
        RECT 1.190 382.520 741.915 385.200 ;
        RECT 4.400 381.120 741.915 382.520 ;
        RECT 1.190 379.120 741.915 381.120 ;
        RECT 4.400 377.720 741.915 379.120 ;
        RECT 1.190 375.040 741.915 377.720 ;
        RECT 4.400 373.640 741.915 375.040 ;
        RECT 1.190 371.640 741.915 373.640 ;
        RECT 4.400 370.240 741.915 371.640 ;
        RECT 1.190 367.560 741.915 370.240 ;
        RECT 4.400 366.160 741.915 367.560 ;
        RECT 1.190 364.160 741.915 366.160 ;
        RECT 4.400 362.760 741.915 364.160 ;
        RECT 1.190 360.080 741.915 362.760 ;
        RECT 4.400 358.680 741.915 360.080 ;
        RECT 1.190 356.680 741.915 358.680 ;
        RECT 4.400 355.280 741.915 356.680 ;
        RECT 1.190 352.600 741.915 355.280 ;
        RECT 4.400 351.200 741.915 352.600 ;
        RECT 1.190 349.200 741.915 351.200 ;
        RECT 4.400 347.800 741.915 349.200 ;
        RECT 1.190 345.120 741.915 347.800 ;
        RECT 4.400 343.720 741.915 345.120 ;
        RECT 1.190 341.720 741.915 343.720 ;
        RECT 4.400 340.320 741.915 341.720 ;
        RECT 1.190 337.640 741.915 340.320 ;
        RECT 4.400 336.240 741.915 337.640 ;
        RECT 1.190 334.240 741.915 336.240 ;
        RECT 4.400 332.840 741.915 334.240 ;
        RECT 1.190 330.160 741.915 332.840 ;
        RECT 4.400 328.760 741.915 330.160 ;
        RECT 1.190 326.760 741.915 328.760 ;
        RECT 4.400 325.360 741.915 326.760 ;
        RECT 1.190 322.680 741.915 325.360 ;
        RECT 4.400 321.280 741.915 322.680 ;
        RECT 1.190 319.280 741.915 321.280 ;
        RECT 4.400 317.880 741.915 319.280 ;
        RECT 1.190 315.200 741.915 317.880 ;
        RECT 4.400 313.800 741.915 315.200 ;
        RECT 1.190 311.800 741.915 313.800 ;
        RECT 4.400 310.400 741.915 311.800 ;
        RECT 1.190 307.720 741.915 310.400 ;
        RECT 4.400 306.320 741.915 307.720 ;
        RECT 1.190 304.320 741.915 306.320 ;
        RECT 4.400 302.920 741.915 304.320 ;
        RECT 1.190 300.920 741.915 302.920 ;
        RECT 4.400 299.520 741.915 300.920 ;
        RECT 1.190 296.840 741.915 299.520 ;
        RECT 4.400 295.440 741.915 296.840 ;
        RECT 1.190 293.440 741.915 295.440 ;
        RECT 4.400 292.040 741.915 293.440 ;
        RECT 1.190 289.360 741.915 292.040 ;
        RECT 4.400 287.960 741.915 289.360 ;
        RECT 1.190 285.960 741.915 287.960 ;
        RECT 4.400 284.560 741.915 285.960 ;
        RECT 1.190 281.880 741.915 284.560 ;
        RECT 4.400 280.480 741.915 281.880 ;
        RECT 1.190 278.480 741.915 280.480 ;
        RECT 4.400 277.080 741.915 278.480 ;
        RECT 1.190 274.400 741.915 277.080 ;
        RECT 4.400 273.000 741.915 274.400 ;
        RECT 1.190 271.000 741.915 273.000 ;
        RECT 4.400 269.600 741.915 271.000 ;
        RECT 1.190 266.920 741.915 269.600 ;
        RECT 4.400 265.520 741.915 266.920 ;
        RECT 1.190 263.520 741.915 265.520 ;
        RECT 4.400 262.120 741.915 263.520 ;
        RECT 1.190 259.440 741.915 262.120 ;
        RECT 4.400 258.040 741.915 259.440 ;
        RECT 1.190 256.040 741.915 258.040 ;
        RECT 4.400 254.640 741.915 256.040 ;
        RECT 1.190 251.960 741.915 254.640 ;
        RECT 4.400 250.560 741.915 251.960 ;
        RECT 1.190 248.560 741.915 250.560 ;
        RECT 4.400 247.160 741.915 248.560 ;
        RECT 1.190 244.480 741.915 247.160 ;
        RECT 4.400 243.080 741.915 244.480 ;
        RECT 1.190 241.080 741.915 243.080 ;
        RECT 4.400 239.680 741.915 241.080 ;
        RECT 1.190 237.000 741.915 239.680 ;
        RECT 4.400 235.600 741.915 237.000 ;
        RECT 1.190 233.600 741.915 235.600 ;
        RECT 4.400 232.200 741.915 233.600 ;
        RECT 1.190 229.520 741.915 232.200 ;
        RECT 4.400 228.120 741.915 229.520 ;
        RECT 1.190 226.120 741.915 228.120 ;
        RECT 4.400 224.720 741.915 226.120 ;
        RECT 1.190 222.040 741.915 224.720 ;
        RECT 4.400 220.640 741.915 222.040 ;
        RECT 1.190 218.640 741.915 220.640 ;
        RECT 4.400 217.240 741.915 218.640 ;
        RECT 1.190 214.560 741.915 217.240 ;
        RECT 4.400 213.160 741.915 214.560 ;
        RECT 1.190 211.160 741.915 213.160 ;
        RECT 4.400 209.760 741.915 211.160 ;
        RECT 1.190 207.080 741.915 209.760 ;
        RECT 4.400 205.680 741.915 207.080 ;
        RECT 1.190 203.680 741.915 205.680 ;
        RECT 4.400 202.280 741.915 203.680 ;
        RECT 1.190 199.600 741.915 202.280 ;
        RECT 4.400 198.200 741.915 199.600 ;
        RECT 1.190 196.200 741.915 198.200 ;
        RECT 4.400 194.800 741.915 196.200 ;
        RECT 1.190 192.120 741.915 194.800 ;
        RECT 4.400 190.720 741.915 192.120 ;
        RECT 1.190 188.720 741.915 190.720 ;
        RECT 4.400 187.320 741.915 188.720 ;
        RECT 1.190 184.640 741.915 187.320 ;
        RECT 4.400 183.240 741.915 184.640 ;
        RECT 1.190 181.240 741.915 183.240 ;
        RECT 4.400 179.840 741.915 181.240 ;
        RECT 1.190 177.160 741.915 179.840 ;
        RECT 4.400 175.760 741.915 177.160 ;
        RECT 1.190 173.760 741.915 175.760 ;
        RECT 4.400 172.360 741.915 173.760 ;
        RECT 1.190 169.680 741.915 172.360 ;
        RECT 4.400 168.280 741.915 169.680 ;
        RECT 1.190 166.280 741.915 168.280 ;
        RECT 4.400 164.880 741.915 166.280 ;
        RECT 1.190 162.200 741.915 164.880 ;
        RECT 4.400 160.800 741.915 162.200 ;
        RECT 1.190 158.800 741.915 160.800 ;
        RECT 4.400 157.400 741.915 158.800 ;
        RECT 1.190 154.720 741.915 157.400 ;
        RECT 4.400 153.320 741.915 154.720 ;
        RECT 1.190 151.320 741.915 153.320 ;
        RECT 4.400 149.920 741.915 151.320 ;
        RECT 1.190 147.920 741.915 149.920 ;
        RECT 4.400 146.520 741.915 147.920 ;
        RECT 1.190 143.840 741.915 146.520 ;
        RECT 4.400 142.440 741.915 143.840 ;
        RECT 1.190 140.440 741.915 142.440 ;
        RECT 4.400 139.040 741.915 140.440 ;
        RECT 1.190 136.360 741.915 139.040 ;
        RECT 4.400 134.960 741.915 136.360 ;
        RECT 1.190 132.960 741.915 134.960 ;
        RECT 4.400 131.560 741.915 132.960 ;
        RECT 1.190 128.880 741.915 131.560 ;
        RECT 4.400 127.480 741.915 128.880 ;
        RECT 1.190 125.480 741.915 127.480 ;
        RECT 4.400 124.080 741.915 125.480 ;
        RECT 1.190 121.400 741.915 124.080 ;
        RECT 4.400 120.000 741.915 121.400 ;
        RECT 1.190 118.000 741.915 120.000 ;
        RECT 4.400 116.600 741.915 118.000 ;
        RECT 1.190 113.920 741.915 116.600 ;
        RECT 4.400 112.520 741.915 113.920 ;
        RECT 1.190 110.520 741.915 112.520 ;
        RECT 4.400 109.120 741.915 110.520 ;
        RECT 1.190 106.440 741.915 109.120 ;
        RECT 4.400 105.040 741.915 106.440 ;
        RECT 1.190 103.040 741.915 105.040 ;
        RECT 4.400 101.640 741.915 103.040 ;
        RECT 1.190 98.960 741.915 101.640 ;
        RECT 4.400 97.560 741.915 98.960 ;
        RECT 1.190 95.560 741.915 97.560 ;
        RECT 4.400 94.160 741.915 95.560 ;
        RECT 1.190 91.480 741.915 94.160 ;
        RECT 4.400 90.080 741.915 91.480 ;
        RECT 1.190 88.080 741.915 90.080 ;
        RECT 4.400 86.680 741.915 88.080 ;
        RECT 1.190 84.000 741.915 86.680 ;
        RECT 4.400 82.600 741.915 84.000 ;
        RECT 1.190 80.600 741.915 82.600 ;
        RECT 4.400 79.200 741.915 80.600 ;
        RECT 1.190 76.520 741.915 79.200 ;
        RECT 4.400 75.120 741.915 76.520 ;
        RECT 1.190 73.120 741.915 75.120 ;
        RECT 4.400 71.720 741.915 73.120 ;
        RECT 1.190 69.040 741.915 71.720 ;
        RECT 4.400 67.640 741.915 69.040 ;
        RECT 1.190 65.640 741.915 67.640 ;
        RECT 4.400 64.240 741.915 65.640 ;
        RECT 1.190 61.560 741.915 64.240 ;
        RECT 4.400 60.160 741.915 61.560 ;
        RECT 1.190 58.160 741.915 60.160 ;
        RECT 4.400 56.760 741.915 58.160 ;
        RECT 1.190 54.080 741.915 56.760 ;
        RECT 4.400 52.680 741.915 54.080 ;
        RECT 1.190 50.680 741.915 52.680 ;
        RECT 4.400 49.280 741.915 50.680 ;
        RECT 1.190 46.600 741.915 49.280 ;
        RECT 4.400 45.200 741.915 46.600 ;
        RECT 1.190 43.200 741.915 45.200 ;
        RECT 4.400 41.800 741.915 43.200 ;
        RECT 1.190 39.120 741.915 41.800 ;
        RECT 4.400 37.720 741.915 39.120 ;
        RECT 1.190 35.720 741.915 37.720 ;
        RECT 4.400 34.320 741.915 35.720 ;
        RECT 1.190 31.640 741.915 34.320 ;
        RECT 4.400 30.240 741.915 31.640 ;
        RECT 1.190 28.240 741.915 30.240 ;
        RECT 4.400 26.840 741.915 28.240 ;
        RECT 1.190 24.160 741.915 26.840 ;
        RECT 4.400 22.760 741.915 24.160 ;
        RECT 1.190 20.760 741.915 22.760 ;
        RECT 4.400 19.360 741.915 20.760 ;
        RECT 1.190 16.680 741.915 19.360 ;
        RECT 4.400 15.280 741.915 16.680 ;
        RECT 1.190 13.280 741.915 15.280 ;
        RECT 4.400 11.880 741.915 13.280 ;
        RECT 1.190 9.200 741.915 11.880 ;
        RECT 4.400 7.800 741.915 9.200 ;
        RECT 1.190 5.800 741.915 7.800 ;
        RECT 4.400 4.400 741.915 5.800 ;
        RECT 1.190 2.400 741.915 4.400 ;
        RECT 4.400 1.535 741.915 2.400 ;
      LAYER met4 ;
        RECT 1.215 737.760 732.945 738.985 ;
        RECT 1.215 10.240 20.640 737.760 ;
        RECT 23.040 10.240 97.440 737.760 ;
        RECT 99.840 10.240 174.240 737.760 ;
        RECT 176.640 10.240 251.040 737.760 ;
        RECT 253.440 10.240 327.840 737.760 ;
        RECT 330.240 10.240 404.640 737.760 ;
        RECT 407.040 10.240 481.440 737.760 ;
        RECT 483.840 10.240 558.240 737.760 ;
        RECT 560.640 10.240 635.040 737.760 ;
        RECT 637.440 10.240 711.840 737.760 ;
        RECT 714.240 10.240 732.945 737.760 ;
        RECT 1.215 6.295 732.945 10.240 ;
  END
END dcache
END LIBRARY

