magic
tech sky130A
magscale 1 2
timestamp 1611821080
<< obsli1 >>
rect 1104 2159 218868 217617
<< obsm1 >>
rect 1104 2128 219498 219632
<< metal2 >>
rect 386 219200 442 220000
rect 1214 219200 1270 220000
rect 2042 219200 2098 220000
rect 2870 219200 2926 220000
rect 3698 219200 3754 220000
rect 4526 219200 4582 220000
rect 5446 219200 5502 220000
rect 6274 219200 6330 220000
rect 7102 219200 7158 220000
rect 7930 219200 7986 220000
rect 8758 219200 8814 220000
rect 9678 219200 9734 220000
rect 10506 219200 10562 220000
rect 11334 219200 11390 220000
rect 12162 219200 12218 220000
rect 12990 219200 13046 220000
rect 13910 219200 13966 220000
rect 14738 219200 14794 220000
rect 15566 219200 15622 220000
rect 16394 219200 16450 220000
rect 17222 219200 17278 220000
rect 18142 219200 18198 220000
rect 18970 219200 19026 220000
rect 19798 219200 19854 220000
rect 20626 219200 20682 220000
rect 21454 219200 21510 220000
rect 22374 219200 22430 220000
rect 23202 219200 23258 220000
rect 24030 219200 24086 220000
rect 24858 219200 24914 220000
rect 25686 219200 25742 220000
rect 26606 219200 26662 220000
rect 27434 219200 27490 220000
rect 28262 219200 28318 220000
rect 29090 219200 29146 220000
rect 29918 219200 29974 220000
rect 30838 219200 30894 220000
rect 31666 219200 31722 220000
rect 32494 219200 32550 220000
rect 33322 219200 33378 220000
rect 34150 219200 34206 220000
rect 35070 219200 35126 220000
rect 35898 219200 35954 220000
rect 36726 219200 36782 220000
rect 37554 219200 37610 220000
rect 38382 219200 38438 220000
rect 39302 219200 39358 220000
rect 40130 219200 40186 220000
rect 40958 219200 41014 220000
rect 41786 219200 41842 220000
rect 42614 219200 42670 220000
rect 43534 219200 43590 220000
rect 44362 219200 44418 220000
rect 45190 219200 45246 220000
rect 46018 219200 46074 220000
rect 46846 219200 46902 220000
rect 47674 219200 47730 220000
rect 48594 219200 48650 220000
rect 49422 219200 49478 220000
rect 50250 219200 50306 220000
rect 51078 219200 51134 220000
rect 51906 219200 51962 220000
rect 52826 219200 52882 220000
rect 53654 219200 53710 220000
rect 54482 219200 54538 220000
rect 55310 219200 55366 220000
rect 56138 219200 56194 220000
rect 57058 219200 57114 220000
rect 57886 219200 57942 220000
rect 58714 219200 58770 220000
rect 59542 219200 59598 220000
rect 60370 219200 60426 220000
rect 61290 219200 61346 220000
rect 62118 219200 62174 220000
rect 62946 219200 63002 220000
rect 63774 219200 63830 220000
rect 64602 219200 64658 220000
rect 65522 219200 65578 220000
rect 66350 219200 66406 220000
rect 67178 219200 67234 220000
rect 68006 219200 68062 220000
rect 68834 219200 68890 220000
rect 69754 219200 69810 220000
rect 70582 219200 70638 220000
rect 71410 219200 71466 220000
rect 72238 219200 72294 220000
rect 73066 219200 73122 220000
rect 73986 219200 74042 220000
rect 74814 219200 74870 220000
rect 75642 219200 75698 220000
rect 76470 219200 76526 220000
rect 77298 219200 77354 220000
rect 78218 219200 78274 220000
rect 79046 219200 79102 220000
rect 79874 219200 79930 220000
rect 80702 219200 80758 220000
rect 81530 219200 81586 220000
rect 82450 219200 82506 220000
rect 83278 219200 83334 220000
rect 84106 219200 84162 220000
rect 84934 219200 84990 220000
rect 85762 219200 85818 220000
rect 86682 219200 86738 220000
rect 87510 219200 87566 220000
rect 88338 219200 88394 220000
rect 89166 219200 89222 220000
rect 89994 219200 90050 220000
rect 90822 219200 90878 220000
rect 91742 219200 91798 220000
rect 92570 219200 92626 220000
rect 93398 219200 93454 220000
rect 94226 219200 94282 220000
rect 95054 219200 95110 220000
rect 95974 219200 96030 220000
rect 96802 219200 96858 220000
rect 97630 219200 97686 220000
rect 98458 219200 98514 220000
rect 99286 219200 99342 220000
rect 100206 219200 100262 220000
rect 101034 219200 101090 220000
rect 101862 219200 101918 220000
rect 102690 219200 102746 220000
rect 103518 219200 103574 220000
rect 104438 219200 104494 220000
rect 105266 219200 105322 220000
rect 106094 219200 106150 220000
rect 106922 219200 106978 220000
rect 107750 219200 107806 220000
rect 108670 219200 108726 220000
rect 109498 219200 109554 220000
rect 110326 219200 110382 220000
rect 111154 219200 111210 220000
rect 111982 219200 112038 220000
rect 112902 219200 112958 220000
rect 113730 219200 113786 220000
rect 114558 219200 114614 220000
rect 115386 219200 115442 220000
rect 116214 219200 116270 220000
rect 117134 219200 117190 220000
rect 117962 219200 118018 220000
rect 118790 219200 118846 220000
rect 119618 219200 119674 220000
rect 120446 219200 120502 220000
rect 121366 219200 121422 220000
rect 122194 219200 122250 220000
rect 123022 219200 123078 220000
rect 123850 219200 123906 220000
rect 124678 219200 124734 220000
rect 125598 219200 125654 220000
rect 126426 219200 126482 220000
rect 127254 219200 127310 220000
rect 128082 219200 128138 220000
rect 128910 219200 128966 220000
rect 129830 219200 129886 220000
rect 130658 219200 130714 220000
rect 131486 219200 131542 220000
rect 132314 219200 132370 220000
rect 133142 219200 133198 220000
rect 133970 219200 134026 220000
rect 134890 219200 134946 220000
rect 135718 219200 135774 220000
rect 136546 219200 136602 220000
rect 137374 219200 137430 220000
rect 138202 219200 138258 220000
rect 139122 219200 139178 220000
rect 139950 219200 140006 220000
rect 140778 219200 140834 220000
rect 141606 219200 141662 220000
rect 142434 219200 142490 220000
rect 143354 219200 143410 220000
rect 144182 219200 144238 220000
rect 145010 219200 145066 220000
rect 145838 219200 145894 220000
rect 146666 219200 146722 220000
rect 147586 219200 147642 220000
rect 148414 219200 148470 220000
rect 149242 219200 149298 220000
rect 150070 219200 150126 220000
rect 150898 219200 150954 220000
rect 151818 219200 151874 220000
rect 152646 219200 152702 220000
rect 153474 219200 153530 220000
rect 154302 219200 154358 220000
rect 155130 219200 155186 220000
rect 156050 219200 156106 220000
rect 156878 219200 156934 220000
rect 157706 219200 157762 220000
rect 158534 219200 158590 220000
rect 159362 219200 159418 220000
rect 160282 219200 160338 220000
rect 161110 219200 161166 220000
rect 161938 219200 161994 220000
rect 162766 219200 162822 220000
rect 163594 219200 163650 220000
rect 164514 219200 164570 220000
rect 165342 219200 165398 220000
rect 166170 219200 166226 220000
rect 166998 219200 167054 220000
rect 167826 219200 167882 220000
rect 168746 219200 168802 220000
rect 169574 219200 169630 220000
rect 170402 219200 170458 220000
rect 171230 219200 171286 220000
rect 172058 219200 172114 220000
rect 172978 219200 173034 220000
rect 173806 219200 173862 220000
rect 174634 219200 174690 220000
rect 175462 219200 175518 220000
rect 176290 219200 176346 220000
rect 177118 219200 177174 220000
rect 178038 219200 178094 220000
rect 178866 219200 178922 220000
rect 179694 219200 179750 220000
rect 180522 219200 180578 220000
rect 181350 219200 181406 220000
rect 182270 219200 182326 220000
rect 183098 219200 183154 220000
rect 183926 219200 183982 220000
rect 184754 219200 184810 220000
rect 185582 219200 185638 220000
rect 186502 219200 186558 220000
rect 187330 219200 187386 220000
rect 188158 219200 188214 220000
rect 188986 219200 189042 220000
rect 189814 219200 189870 220000
rect 190734 219200 190790 220000
rect 191562 219200 191618 220000
rect 192390 219200 192446 220000
rect 193218 219200 193274 220000
rect 194046 219200 194102 220000
rect 194966 219200 195022 220000
rect 195794 219200 195850 220000
rect 196622 219200 196678 220000
rect 197450 219200 197506 220000
rect 198278 219200 198334 220000
rect 199198 219200 199254 220000
rect 200026 219200 200082 220000
rect 200854 219200 200910 220000
rect 201682 219200 201738 220000
rect 202510 219200 202566 220000
rect 203430 219200 203486 220000
rect 204258 219200 204314 220000
rect 205086 219200 205142 220000
rect 205914 219200 205970 220000
rect 206742 219200 206798 220000
rect 207662 219200 207718 220000
rect 208490 219200 208546 220000
rect 209318 219200 209374 220000
rect 210146 219200 210202 220000
rect 210974 219200 211030 220000
rect 211894 219200 211950 220000
rect 212722 219200 212778 220000
rect 213550 219200 213606 220000
rect 214378 219200 214434 220000
rect 215206 219200 215262 220000
rect 216126 219200 216182 220000
rect 216954 219200 217010 220000
rect 217782 219200 217838 220000
rect 218610 219200 218666 220000
rect 219438 219200 219494 220000
<< obsm2 >>
rect 18 219144 330 219638
rect 498 219144 1158 219638
rect 1326 219144 1986 219638
rect 2154 219144 2814 219638
rect 2982 219144 3642 219638
rect 3810 219144 4470 219638
rect 4638 219144 5390 219638
rect 5558 219144 6218 219638
rect 6386 219144 7046 219638
rect 7214 219144 7874 219638
rect 8042 219144 8702 219638
rect 8870 219144 9622 219638
rect 9790 219144 10450 219638
rect 10618 219144 11278 219638
rect 11446 219144 12106 219638
rect 12274 219144 12934 219638
rect 13102 219144 13854 219638
rect 14022 219144 14682 219638
rect 14850 219144 15510 219638
rect 15678 219144 16338 219638
rect 16506 219144 17166 219638
rect 17334 219144 18086 219638
rect 18254 219144 18914 219638
rect 19082 219144 19742 219638
rect 19910 219144 20570 219638
rect 20738 219144 21398 219638
rect 21566 219144 22318 219638
rect 22486 219144 23146 219638
rect 23314 219144 23974 219638
rect 24142 219144 24802 219638
rect 24970 219144 25630 219638
rect 25798 219144 26550 219638
rect 26718 219144 27378 219638
rect 27546 219144 28206 219638
rect 28374 219144 29034 219638
rect 29202 219144 29862 219638
rect 30030 219144 30782 219638
rect 30950 219144 31610 219638
rect 31778 219144 32438 219638
rect 32606 219144 33266 219638
rect 33434 219144 34094 219638
rect 34262 219144 35014 219638
rect 35182 219144 35842 219638
rect 36010 219144 36670 219638
rect 36838 219144 37498 219638
rect 37666 219144 38326 219638
rect 38494 219144 39246 219638
rect 39414 219144 40074 219638
rect 40242 219144 40902 219638
rect 41070 219144 41730 219638
rect 41898 219144 42558 219638
rect 42726 219144 43478 219638
rect 43646 219144 44306 219638
rect 44474 219144 45134 219638
rect 45302 219144 45962 219638
rect 46130 219144 46790 219638
rect 46958 219144 47618 219638
rect 47786 219144 48538 219638
rect 48706 219144 49366 219638
rect 49534 219144 50194 219638
rect 50362 219144 51022 219638
rect 51190 219144 51850 219638
rect 52018 219144 52770 219638
rect 52938 219144 53598 219638
rect 53766 219144 54426 219638
rect 54594 219144 55254 219638
rect 55422 219144 56082 219638
rect 56250 219144 57002 219638
rect 57170 219144 57830 219638
rect 57998 219144 58658 219638
rect 58826 219144 59486 219638
rect 59654 219144 60314 219638
rect 60482 219144 61234 219638
rect 61402 219144 62062 219638
rect 62230 219144 62890 219638
rect 63058 219144 63718 219638
rect 63886 219144 64546 219638
rect 64714 219144 65466 219638
rect 65634 219144 66294 219638
rect 66462 219144 67122 219638
rect 67290 219144 67950 219638
rect 68118 219144 68778 219638
rect 68946 219144 69698 219638
rect 69866 219144 70526 219638
rect 70694 219144 71354 219638
rect 71522 219144 72182 219638
rect 72350 219144 73010 219638
rect 73178 219144 73930 219638
rect 74098 219144 74758 219638
rect 74926 219144 75586 219638
rect 75754 219144 76414 219638
rect 76582 219144 77242 219638
rect 77410 219144 78162 219638
rect 78330 219144 78990 219638
rect 79158 219144 79818 219638
rect 79986 219144 80646 219638
rect 80814 219144 81474 219638
rect 81642 219144 82394 219638
rect 82562 219144 83222 219638
rect 83390 219144 84050 219638
rect 84218 219144 84878 219638
rect 85046 219144 85706 219638
rect 85874 219144 86626 219638
rect 86794 219144 87454 219638
rect 87622 219144 88282 219638
rect 88450 219144 89110 219638
rect 89278 219144 89938 219638
rect 90106 219144 90766 219638
rect 90934 219144 91686 219638
rect 91854 219144 92514 219638
rect 92682 219144 93342 219638
rect 93510 219144 94170 219638
rect 94338 219144 94998 219638
rect 95166 219144 95918 219638
rect 96086 219144 96746 219638
rect 96914 219144 97574 219638
rect 97742 219144 98402 219638
rect 98570 219144 99230 219638
rect 99398 219144 100150 219638
rect 100318 219144 100978 219638
rect 101146 219144 101806 219638
rect 101974 219144 102634 219638
rect 102802 219144 103462 219638
rect 103630 219144 104382 219638
rect 104550 219144 105210 219638
rect 105378 219144 106038 219638
rect 106206 219144 106866 219638
rect 107034 219144 107694 219638
rect 107862 219144 108614 219638
rect 108782 219144 109442 219638
rect 109610 219144 110270 219638
rect 110438 219144 111098 219638
rect 111266 219144 111926 219638
rect 112094 219144 112846 219638
rect 113014 219144 113674 219638
rect 113842 219144 114502 219638
rect 114670 219144 115330 219638
rect 115498 219144 116158 219638
rect 116326 219144 117078 219638
rect 117246 219144 117906 219638
rect 118074 219144 118734 219638
rect 118902 219144 119562 219638
rect 119730 219144 120390 219638
rect 120558 219144 121310 219638
rect 121478 219144 122138 219638
rect 122306 219144 122966 219638
rect 123134 219144 123794 219638
rect 123962 219144 124622 219638
rect 124790 219144 125542 219638
rect 125710 219144 126370 219638
rect 126538 219144 127198 219638
rect 127366 219144 128026 219638
rect 128194 219144 128854 219638
rect 129022 219144 129774 219638
rect 129942 219144 130602 219638
rect 130770 219144 131430 219638
rect 131598 219144 132258 219638
rect 132426 219144 133086 219638
rect 133254 219144 133914 219638
rect 134082 219144 134834 219638
rect 135002 219144 135662 219638
rect 135830 219144 136490 219638
rect 136658 219144 137318 219638
rect 137486 219144 138146 219638
rect 138314 219144 139066 219638
rect 139234 219144 139894 219638
rect 140062 219144 140722 219638
rect 140890 219144 141550 219638
rect 141718 219144 142378 219638
rect 142546 219144 143298 219638
rect 143466 219144 144126 219638
rect 144294 219144 144954 219638
rect 145122 219144 145782 219638
rect 145950 219144 146610 219638
rect 146778 219144 147530 219638
rect 147698 219144 148358 219638
rect 148526 219144 149186 219638
rect 149354 219144 150014 219638
rect 150182 219144 150842 219638
rect 151010 219144 151762 219638
rect 151930 219144 152590 219638
rect 152758 219144 153418 219638
rect 153586 219144 154246 219638
rect 154414 219144 155074 219638
rect 155242 219144 155994 219638
rect 156162 219144 156822 219638
rect 156990 219144 157650 219638
rect 157818 219144 158478 219638
rect 158646 219144 159306 219638
rect 159474 219144 160226 219638
rect 160394 219144 161054 219638
rect 161222 219144 161882 219638
rect 162050 219144 162710 219638
rect 162878 219144 163538 219638
rect 163706 219144 164458 219638
rect 164626 219144 165286 219638
rect 165454 219144 166114 219638
rect 166282 219144 166942 219638
rect 167110 219144 167770 219638
rect 167938 219144 168690 219638
rect 168858 219144 169518 219638
rect 169686 219144 170346 219638
rect 170514 219144 171174 219638
rect 171342 219144 172002 219638
rect 172170 219144 172922 219638
rect 173090 219144 173750 219638
rect 173918 219144 174578 219638
rect 174746 219144 175406 219638
rect 175574 219144 176234 219638
rect 176402 219144 177062 219638
rect 177230 219144 177982 219638
rect 178150 219144 178810 219638
rect 178978 219144 179638 219638
rect 179806 219144 180466 219638
rect 180634 219144 181294 219638
rect 181462 219144 182214 219638
rect 182382 219144 183042 219638
rect 183210 219144 183870 219638
rect 184038 219144 184698 219638
rect 184866 219144 185526 219638
rect 185694 219144 186446 219638
rect 186614 219144 187274 219638
rect 187442 219144 188102 219638
rect 188270 219144 188930 219638
rect 189098 219144 189758 219638
rect 189926 219144 190678 219638
rect 190846 219144 191506 219638
rect 191674 219144 192334 219638
rect 192502 219144 193162 219638
rect 193330 219144 193990 219638
rect 194158 219144 194910 219638
rect 195078 219144 195738 219638
rect 195906 219144 196566 219638
rect 196734 219144 197394 219638
rect 197562 219144 198222 219638
rect 198390 219144 199142 219638
rect 199310 219144 199970 219638
rect 200138 219144 200798 219638
rect 200966 219144 201626 219638
rect 201794 219144 202454 219638
rect 202622 219144 203374 219638
rect 203542 219144 204202 219638
rect 204370 219144 205030 219638
rect 205198 219144 205858 219638
rect 206026 219144 206686 219638
rect 206854 219144 207606 219638
rect 207774 219144 208434 219638
rect 208602 219144 209262 219638
rect 209430 219144 210090 219638
rect 210258 219144 210918 219638
rect 211086 219144 211838 219638
rect 212006 219144 212666 219638
rect 212834 219144 213494 219638
rect 213662 219144 214322 219638
rect 214490 219144 215150 219638
rect 215318 219144 216070 219638
rect 216238 219144 216898 219638
rect 217066 219144 217726 219638
rect 217894 219144 218554 219638
rect 218722 219144 219382 219638
rect 18 847 219492 219144
<< metal3 >>
rect 219200 219104 220000 219224
rect 219200 217472 220000 217592
rect 219200 215704 220000 215824
rect 219200 214072 220000 214192
rect 219200 212304 220000 212424
rect 219200 210672 220000 210792
rect 219200 208904 220000 209024
rect 219200 207272 220000 207392
rect 219200 205504 220000 205624
rect 219200 203872 220000 203992
rect 219200 202240 220000 202360
rect 219200 200472 220000 200592
rect 219200 198840 220000 198960
rect 219200 197072 220000 197192
rect 219200 195440 220000 195560
rect 219200 193672 220000 193792
rect 219200 192040 220000 192160
rect 219200 190272 220000 190392
rect 219200 188640 220000 188760
rect 219200 187008 220000 187128
rect 219200 185240 220000 185360
rect 219200 183608 220000 183728
rect 219200 181840 220000 181960
rect 219200 180208 220000 180328
rect 219200 178440 220000 178560
rect 219200 176808 220000 176928
rect 219200 175040 220000 175160
rect 219200 173408 220000 173528
rect 219200 171776 220000 171896
rect 219200 170008 220000 170128
rect 219200 168376 220000 168496
rect 219200 166608 220000 166728
rect 219200 164976 220000 165096
rect 219200 163208 220000 163328
rect 219200 161576 220000 161696
rect 219200 159808 220000 159928
rect 219200 158176 220000 158296
rect 219200 156544 220000 156664
rect 219200 154776 220000 154896
rect 219200 153144 220000 153264
rect 219200 151376 220000 151496
rect 219200 149744 220000 149864
rect 219200 147976 220000 148096
rect 219200 146344 220000 146464
rect 219200 144576 220000 144696
rect 219200 142944 220000 143064
rect 219200 141312 220000 141432
rect 219200 139544 220000 139664
rect 219200 137912 220000 138032
rect 219200 136144 220000 136264
rect 219200 134512 220000 134632
rect 219200 132744 220000 132864
rect 219200 131112 220000 131232
rect 219200 129344 220000 129464
rect 219200 127712 220000 127832
rect 219200 126080 220000 126200
rect 219200 124312 220000 124432
rect 219200 122680 220000 122800
rect 219200 120912 220000 121032
rect 219200 119280 220000 119400
rect 219200 117512 220000 117632
rect 219200 115880 220000 116000
rect 219200 114112 220000 114232
rect 219200 112480 220000 112600
rect 219200 110848 220000 110968
rect 219200 109080 220000 109200
rect 219200 107448 220000 107568
rect 219200 105680 220000 105800
rect 219200 104048 220000 104168
rect 219200 102280 220000 102400
rect 219200 100648 220000 100768
rect 219200 98880 220000 99000
rect 219200 97248 220000 97368
rect 219200 95480 220000 95600
rect 219200 93848 220000 93968
rect 219200 92216 220000 92336
rect 219200 90448 220000 90568
rect 219200 88816 220000 88936
rect 219200 87048 220000 87168
rect 219200 85416 220000 85536
rect 219200 83648 220000 83768
rect 219200 82016 220000 82136
rect 219200 80248 220000 80368
rect 219200 78616 220000 78736
rect 219200 76984 220000 77104
rect 219200 75216 220000 75336
rect 219200 73584 220000 73704
rect 219200 71816 220000 71936
rect 219200 70184 220000 70304
rect 219200 68416 220000 68536
rect 219200 66784 220000 66904
rect 219200 65016 220000 65136
rect 219200 63384 220000 63504
rect 219200 61752 220000 61872
rect 219200 59984 220000 60104
rect 219200 58352 220000 58472
rect 219200 56584 220000 56704
rect 219200 54952 220000 55072
rect 219200 53184 220000 53304
rect 219200 51552 220000 51672
rect 219200 49784 220000 49904
rect 219200 48152 220000 48272
rect 219200 46520 220000 46640
rect 219200 44752 220000 44872
rect 219200 43120 220000 43240
rect 219200 41352 220000 41472
rect 219200 39720 220000 39840
rect 219200 37952 220000 38072
rect 219200 36320 220000 36440
rect 219200 34552 220000 34672
rect 219200 32920 220000 33040
rect 219200 31288 220000 31408
rect 219200 29520 220000 29640
rect 219200 27888 220000 28008
rect 219200 26120 220000 26240
rect 219200 24488 220000 24608
rect 219200 22720 220000 22840
rect 219200 21088 220000 21208
rect 219200 19320 220000 19440
rect 219200 17688 220000 17808
rect 219200 16056 220000 16176
rect 219200 14288 220000 14408
rect 219200 12656 220000 12776
rect 219200 10888 220000 11008
rect 219200 9256 220000 9376
rect 219200 7488 220000 7608
rect 219200 5856 220000 5976
rect 219200 4088 220000 4208
rect 219200 2456 220000 2576
rect 219200 824 220000 944
<< obsm3 >>
rect 13 219024 219120 219197
rect 13 217672 219200 219024
rect 13 217392 219120 217672
rect 13 215904 219200 217392
rect 13 215624 219120 215904
rect 13 214272 219200 215624
rect 13 213992 219120 214272
rect 13 212504 219200 213992
rect 13 212224 219120 212504
rect 13 210872 219200 212224
rect 13 210592 219120 210872
rect 13 209104 219200 210592
rect 13 208824 219120 209104
rect 13 207472 219200 208824
rect 13 207192 219120 207472
rect 13 205704 219200 207192
rect 13 205424 219120 205704
rect 13 204072 219200 205424
rect 13 203792 219120 204072
rect 13 202440 219200 203792
rect 13 202160 219120 202440
rect 13 200672 219200 202160
rect 13 200392 219120 200672
rect 13 199040 219200 200392
rect 13 198760 219120 199040
rect 13 197272 219200 198760
rect 13 196992 219120 197272
rect 13 195640 219200 196992
rect 13 195360 219120 195640
rect 13 193872 219200 195360
rect 13 193592 219120 193872
rect 13 192240 219200 193592
rect 13 191960 219120 192240
rect 13 190472 219200 191960
rect 13 190192 219120 190472
rect 13 188840 219200 190192
rect 13 188560 219120 188840
rect 13 187208 219200 188560
rect 13 186928 219120 187208
rect 13 185440 219200 186928
rect 13 185160 219120 185440
rect 13 183808 219200 185160
rect 13 183528 219120 183808
rect 13 182040 219200 183528
rect 13 181760 219120 182040
rect 13 180408 219200 181760
rect 13 180128 219120 180408
rect 13 178640 219200 180128
rect 13 178360 219120 178640
rect 13 177008 219200 178360
rect 13 176728 219120 177008
rect 13 175240 219200 176728
rect 13 174960 219120 175240
rect 13 173608 219200 174960
rect 13 173328 219120 173608
rect 13 171976 219200 173328
rect 13 171696 219120 171976
rect 13 170208 219200 171696
rect 13 169928 219120 170208
rect 13 168576 219200 169928
rect 13 168296 219120 168576
rect 13 166808 219200 168296
rect 13 166528 219120 166808
rect 13 165176 219200 166528
rect 13 164896 219120 165176
rect 13 163408 219200 164896
rect 13 163128 219120 163408
rect 13 161776 219200 163128
rect 13 161496 219120 161776
rect 13 160008 219200 161496
rect 13 159728 219120 160008
rect 13 158376 219200 159728
rect 13 158096 219120 158376
rect 13 156744 219200 158096
rect 13 156464 219120 156744
rect 13 154976 219200 156464
rect 13 154696 219120 154976
rect 13 153344 219200 154696
rect 13 153064 219120 153344
rect 13 151576 219200 153064
rect 13 151296 219120 151576
rect 13 149944 219200 151296
rect 13 149664 219120 149944
rect 13 148176 219200 149664
rect 13 147896 219120 148176
rect 13 146544 219200 147896
rect 13 146264 219120 146544
rect 13 144776 219200 146264
rect 13 144496 219120 144776
rect 13 143144 219200 144496
rect 13 142864 219120 143144
rect 13 141512 219200 142864
rect 13 141232 219120 141512
rect 13 139744 219200 141232
rect 13 139464 219120 139744
rect 13 138112 219200 139464
rect 13 137832 219120 138112
rect 13 136344 219200 137832
rect 13 136064 219120 136344
rect 13 134712 219200 136064
rect 13 134432 219120 134712
rect 13 132944 219200 134432
rect 13 132664 219120 132944
rect 13 131312 219200 132664
rect 13 131032 219120 131312
rect 13 129544 219200 131032
rect 13 129264 219120 129544
rect 13 127912 219200 129264
rect 13 127632 219120 127912
rect 13 126280 219200 127632
rect 13 126000 219120 126280
rect 13 124512 219200 126000
rect 13 124232 219120 124512
rect 13 122880 219200 124232
rect 13 122600 219120 122880
rect 13 121112 219200 122600
rect 13 120832 219120 121112
rect 13 119480 219200 120832
rect 13 119200 219120 119480
rect 13 117712 219200 119200
rect 13 117432 219120 117712
rect 13 116080 219200 117432
rect 13 115800 219120 116080
rect 13 114312 219200 115800
rect 13 114032 219120 114312
rect 13 112680 219200 114032
rect 13 112400 219120 112680
rect 13 111048 219200 112400
rect 13 110768 219120 111048
rect 13 109280 219200 110768
rect 13 109000 219120 109280
rect 13 107648 219200 109000
rect 13 107368 219120 107648
rect 13 105880 219200 107368
rect 13 105600 219120 105880
rect 13 104248 219200 105600
rect 13 103968 219120 104248
rect 13 102480 219200 103968
rect 13 102200 219120 102480
rect 13 100848 219200 102200
rect 13 100568 219120 100848
rect 13 99080 219200 100568
rect 13 98800 219120 99080
rect 13 97448 219200 98800
rect 13 97168 219120 97448
rect 13 95680 219200 97168
rect 13 95400 219120 95680
rect 13 94048 219200 95400
rect 13 93768 219120 94048
rect 13 92416 219200 93768
rect 13 92136 219120 92416
rect 13 90648 219200 92136
rect 13 90368 219120 90648
rect 13 89016 219200 90368
rect 13 88736 219120 89016
rect 13 87248 219200 88736
rect 13 86968 219120 87248
rect 13 85616 219200 86968
rect 13 85336 219120 85616
rect 13 83848 219200 85336
rect 13 83568 219120 83848
rect 13 82216 219200 83568
rect 13 81936 219120 82216
rect 13 80448 219200 81936
rect 13 80168 219120 80448
rect 13 78816 219200 80168
rect 13 78536 219120 78816
rect 13 77184 219200 78536
rect 13 76904 219120 77184
rect 13 75416 219200 76904
rect 13 75136 219120 75416
rect 13 73784 219200 75136
rect 13 73504 219120 73784
rect 13 72016 219200 73504
rect 13 71736 219120 72016
rect 13 70384 219200 71736
rect 13 70104 219120 70384
rect 13 68616 219200 70104
rect 13 68336 219120 68616
rect 13 66984 219200 68336
rect 13 66704 219120 66984
rect 13 65216 219200 66704
rect 13 64936 219120 65216
rect 13 63584 219200 64936
rect 13 63304 219120 63584
rect 13 61952 219200 63304
rect 13 61672 219120 61952
rect 13 60184 219200 61672
rect 13 59904 219120 60184
rect 13 58552 219200 59904
rect 13 58272 219120 58552
rect 13 56784 219200 58272
rect 13 56504 219120 56784
rect 13 55152 219200 56504
rect 13 54872 219120 55152
rect 13 53384 219200 54872
rect 13 53104 219120 53384
rect 13 51752 219200 53104
rect 13 51472 219120 51752
rect 13 49984 219200 51472
rect 13 49704 219120 49984
rect 13 48352 219200 49704
rect 13 48072 219120 48352
rect 13 46720 219200 48072
rect 13 46440 219120 46720
rect 13 44952 219200 46440
rect 13 44672 219120 44952
rect 13 43320 219200 44672
rect 13 43040 219120 43320
rect 13 41552 219200 43040
rect 13 41272 219120 41552
rect 13 39920 219200 41272
rect 13 39640 219120 39920
rect 13 38152 219200 39640
rect 13 37872 219120 38152
rect 13 36520 219200 37872
rect 13 36240 219120 36520
rect 13 34752 219200 36240
rect 13 34472 219120 34752
rect 13 33120 219200 34472
rect 13 32840 219120 33120
rect 13 31488 219200 32840
rect 13 31208 219120 31488
rect 13 29720 219200 31208
rect 13 29440 219120 29720
rect 13 28088 219200 29440
rect 13 27808 219120 28088
rect 13 26320 219200 27808
rect 13 26040 219120 26320
rect 13 24688 219200 26040
rect 13 24408 219120 24688
rect 13 22920 219200 24408
rect 13 22640 219120 22920
rect 13 21288 219200 22640
rect 13 21008 219120 21288
rect 13 19520 219200 21008
rect 13 19240 219120 19520
rect 13 17888 219200 19240
rect 13 17608 219120 17888
rect 13 16256 219200 17608
rect 13 15976 219120 16256
rect 13 14488 219200 15976
rect 13 14208 219120 14488
rect 13 12856 219200 14208
rect 13 12576 219120 12856
rect 13 11088 219200 12576
rect 13 10808 219120 11088
rect 13 9456 219200 10808
rect 13 9176 219120 9456
rect 13 7688 219200 9176
rect 13 7408 219120 7688
rect 13 6056 219200 7408
rect 13 5776 219120 6056
rect 13 4288 219200 5776
rect 13 4008 219120 4288
rect 13 2656 219200 4008
rect 13 2376 219120 2656
rect 13 1024 219200 2376
rect 13 851 219120 1024
<< metal4 >>
rect 4208 2128 4528 217648
rect 19568 2128 19888 217648
rect 34928 2128 35248 217648
rect 50288 2128 50608 217648
rect 65648 2128 65968 217648
rect 81008 2128 81328 217648
rect 96368 2128 96688 217648
rect 111728 2128 112048 217648
rect 127088 2128 127408 217648
rect 142448 2128 142768 217648
rect 157808 2128 158128 217648
rect 173168 2128 173488 217648
rect 188528 2128 188848 217648
rect 203888 2128 204208 217648
<< obsm4 >>
rect 3555 13771 4128 217157
rect 4608 13771 19488 217157
rect 19968 13771 34848 217157
rect 35328 13771 50208 217157
rect 50688 13771 65568 217157
rect 66048 13771 80928 217157
rect 81408 13771 96288 217157
rect 96768 13771 111648 217157
rect 112128 13771 127008 217157
rect 127488 13771 142368 217157
rect 142848 13771 157728 217157
rect 158208 13771 173088 217157
rect 173568 13771 188448 217157
rect 188928 13771 203808 217157
rect 204288 13771 217981 217157
<< labels >>
rlabel metal2 s 386 219200 442 220000 6 clk
port 1 nsew signal input
rlabel metal2 s 1214 219200 1270 220000 6 m_in[0]
port 2 nsew signal input
rlabel metal2 s 85762 219200 85818 220000 6 m_in[100]
port 3 nsew signal input
rlabel metal2 s 86682 219200 86738 220000 6 m_in[101]
port 4 nsew signal input
rlabel metal2 s 87510 219200 87566 220000 6 m_in[102]
port 5 nsew signal input
rlabel metal2 s 88338 219200 88394 220000 6 m_in[103]
port 6 nsew signal input
rlabel metal2 s 89166 219200 89222 220000 6 m_in[104]
port 7 nsew signal input
rlabel metal2 s 89994 219200 90050 220000 6 m_in[105]
port 8 nsew signal input
rlabel metal2 s 90822 219200 90878 220000 6 m_in[106]
port 9 nsew signal input
rlabel metal2 s 91742 219200 91798 220000 6 m_in[107]
port 10 nsew signal input
rlabel metal2 s 92570 219200 92626 220000 6 m_in[108]
port 11 nsew signal input
rlabel metal2 s 93398 219200 93454 220000 6 m_in[109]
port 12 nsew signal input
rlabel metal2 s 9678 219200 9734 220000 6 m_in[10]
port 13 nsew signal input
rlabel metal2 s 94226 219200 94282 220000 6 m_in[110]
port 14 nsew signal input
rlabel metal2 s 95054 219200 95110 220000 6 m_in[111]
port 15 nsew signal input
rlabel metal2 s 95974 219200 96030 220000 6 m_in[112]
port 16 nsew signal input
rlabel metal2 s 96802 219200 96858 220000 6 m_in[113]
port 17 nsew signal input
rlabel metal2 s 97630 219200 97686 220000 6 m_in[114]
port 18 nsew signal input
rlabel metal2 s 98458 219200 98514 220000 6 m_in[115]
port 19 nsew signal input
rlabel metal2 s 99286 219200 99342 220000 6 m_in[116]
port 20 nsew signal input
rlabel metal2 s 100206 219200 100262 220000 6 m_in[117]
port 21 nsew signal input
rlabel metal2 s 101034 219200 101090 220000 6 m_in[118]
port 22 nsew signal input
rlabel metal2 s 101862 219200 101918 220000 6 m_in[119]
port 23 nsew signal input
rlabel metal2 s 10506 219200 10562 220000 6 m_in[11]
port 24 nsew signal input
rlabel metal2 s 102690 219200 102746 220000 6 m_in[120]
port 25 nsew signal input
rlabel metal2 s 103518 219200 103574 220000 6 m_in[121]
port 26 nsew signal input
rlabel metal2 s 104438 219200 104494 220000 6 m_in[122]
port 27 nsew signal input
rlabel metal2 s 105266 219200 105322 220000 6 m_in[123]
port 28 nsew signal input
rlabel metal2 s 106094 219200 106150 220000 6 m_in[124]
port 29 nsew signal input
rlabel metal2 s 106922 219200 106978 220000 6 m_in[125]
port 30 nsew signal input
rlabel metal2 s 107750 219200 107806 220000 6 m_in[126]
port 31 nsew signal input
rlabel metal2 s 108670 219200 108726 220000 6 m_in[127]
port 32 nsew signal input
rlabel metal2 s 109498 219200 109554 220000 6 m_in[128]
port 33 nsew signal input
rlabel metal2 s 110326 219200 110382 220000 6 m_in[129]
port 34 nsew signal input
rlabel metal2 s 11334 219200 11390 220000 6 m_in[12]
port 35 nsew signal input
rlabel metal2 s 111154 219200 111210 220000 6 m_in[130]
port 36 nsew signal input
rlabel metal2 s 111982 219200 112038 220000 6 m_in[131]
port 37 nsew signal input
rlabel metal2 s 112902 219200 112958 220000 6 m_in[132]
port 38 nsew signal input
rlabel metal2 s 113730 219200 113786 220000 6 m_in[133]
port 39 nsew signal input
rlabel metal2 s 114558 219200 114614 220000 6 m_in[134]
port 40 nsew signal input
rlabel metal2 s 115386 219200 115442 220000 6 m_in[135]
port 41 nsew signal input
rlabel metal2 s 116214 219200 116270 220000 6 m_in[136]
port 42 nsew signal input
rlabel metal2 s 117134 219200 117190 220000 6 m_in[137]
port 43 nsew signal input
rlabel metal2 s 117962 219200 118018 220000 6 m_in[138]
port 44 nsew signal input
rlabel metal2 s 118790 219200 118846 220000 6 m_in[139]
port 45 nsew signal input
rlabel metal2 s 12162 219200 12218 220000 6 m_in[13]
port 46 nsew signal input
rlabel metal2 s 119618 219200 119674 220000 6 m_in[140]
port 47 nsew signal input
rlabel metal2 s 120446 219200 120502 220000 6 m_in[141]
port 48 nsew signal input
rlabel metal2 s 121366 219200 121422 220000 6 m_in[142]
port 49 nsew signal input
rlabel metal2 s 122194 219200 122250 220000 6 m_in[143]
port 50 nsew signal input
rlabel metal2 s 123022 219200 123078 220000 6 m_in[144]
port 51 nsew signal input
rlabel metal2 s 123850 219200 123906 220000 6 m_in[145]
port 52 nsew signal input
rlabel metal2 s 124678 219200 124734 220000 6 m_in[146]
port 53 nsew signal input
rlabel metal2 s 125598 219200 125654 220000 6 m_in[147]
port 54 nsew signal input
rlabel metal2 s 126426 219200 126482 220000 6 m_in[148]
port 55 nsew signal input
rlabel metal2 s 127254 219200 127310 220000 6 m_in[149]
port 56 nsew signal input
rlabel metal2 s 12990 219200 13046 220000 6 m_in[14]
port 57 nsew signal input
rlabel metal2 s 128082 219200 128138 220000 6 m_in[150]
port 58 nsew signal input
rlabel metal2 s 128910 219200 128966 220000 6 m_in[151]
port 59 nsew signal input
rlabel metal2 s 129830 219200 129886 220000 6 m_in[152]
port 60 nsew signal input
rlabel metal2 s 130658 219200 130714 220000 6 m_in[153]
port 61 nsew signal input
rlabel metal2 s 131486 219200 131542 220000 6 m_in[154]
port 62 nsew signal input
rlabel metal2 s 132314 219200 132370 220000 6 m_in[155]
port 63 nsew signal input
rlabel metal2 s 133142 219200 133198 220000 6 m_in[156]
port 64 nsew signal input
rlabel metal2 s 133970 219200 134026 220000 6 m_in[157]
port 65 nsew signal input
rlabel metal2 s 134890 219200 134946 220000 6 m_in[158]
port 66 nsew signal input
rlabel metal2 s 135718 219200 135774 220000 6 m_in[159]
port 67 nsew signal input
rlabel metal2 s 13910 219200 13966 220000 6 m_in[15]
port 68 nsew signal input
rlabel metal2 s 136546 219200 136602 220000 6 m_in[160]
port 69 nsew signal input
rlabel metal2 s 137374 219200 137430 220000 6 m_in[161]
port 70 nsew signal input
rlabel metal2 s 138202 219200 138258 220000 6 m_in[162]
port 71 nsew signal input
rlabel metal2 s 139122 219200 139178 220000 6 m_in[163]
port 72 nsew signal input
rlabel metal2 s 139950 219200 140006 220000 6 m_in[164]
port 73 nsew signal input
rlabel metal2 s 140778 219200 140834 220000 6 m_in[165]
port 74 nsew signal input
rlabel metal2 s 141606 219200 141662 220000 6 m_in[166]
port 75 nsew signal input
rlabel metal2 s 142434 219200 142490 220000 6 m_in[167]
port 76 nsew signal input
rlabel metal2 s 143354 219200 143410 220000 6 m_in[168]
port 77 nsew signal input
rlabel metal2 s 144182 219200 144238 220000 6 m_in[169]
port 78 nsew signal input
rlabel metal2 s 14738 219200 14794 220000 6 m_in[16]
port 79 nsew signal input
rlabel metal2 s 145010 219200 145066 220000 6 m_in[170]
port 80 nsew signal input
rlabel metal2 s 145838 219200 145894 220000 6 m_in[171]
port 81 nsew signal input
rlabel metal2 s 146666 219200 146722 220000 6 m_in[172]
port 82 nsew signal input
rlabel metal2 s 147586 219200 147642 220000 6 m_in[173]
port 83 nsew signal input
rlabel metal2 s 148414 219200 148470 220000 6 m_in[174]
port 84 nsew signal input
rlabel metal2 s 149242 219200 149298 220000 6 m_in[175]
port 85 nsew signal input
rlabel metal2 s 150070 219200 150126 220000 6 m_in[176]
port 86 nsew signal input
rlabel metal2 s 150898 219200 150954 220000 6 m_in[177]
port 87 nsew signal input
rlabel metal2 s 151818 219200 151874 220000 6 m_in[178]
port 88 nsew signal input
rlabel metal2 s 152646 219200 152702 220000 6 m_in[179]
port 89 nsew signal input
rlabel metal2 s 15566 219200 15622 220000 6 m_in[17]
port 90 nsew signal input
rlabel metal2 s 153474 219200 153530 220000 6 m_in[180]
port 91 nsew signal input
rlabel metal2 s 154302 219200 154358 220000 6 m_in[181]
port 92 nsew signal input
rlabel metal2 s 155130 219200 155186 220000 6 m_in[182]
port 93 nsew signal input
rlabel metal2 s 156050 219200 156106 220000 6 m_in[183]
port 94 nsew signal input
rlabel metal2 s 156878 219200 156934 220000 6 m_in[184]
port 95 nsew signal input
rlabel metal2 s 157706 219200 157762 220000 6 m_in[185]
port 96 nsew signal input
rlabel metal2 s 158534 219200 158590 220000 6 m_in[186]
port 97 nsew signal input
rlabel metal2 s 159362 219200 159418 220000 6 m_in[187]
port 98 nsew signal input
rlabel metal2 s 160282 219200 160338 220000 6 m_in[188]
port 99 nsew signal input
rlabel metal2 s 161110 219200 161166 220000 6 m_in[189]
port 100 nsew signal input
rlabel metal2 s 16394 219200 16450 220000 6 m_in[18]
port 101 nsew signal input
rlabel metal2 s 161938 219200 161994 220000 6 m_in[190]
port 102 nsew signal input
rlabel metal2 s 162766 219200 162822 220000 6 m_in[191]
port 103 nsew signal input
rlabel metal2 s 163594 219200 163650 220000 6 m_in[192]
port 104 nsew signal input
rlabel metal2 s 164514 219200 164570 220000 6 m_in[193]
port 105 nsew signal input
rlabel metal2 s 165342 219200 165398 220000 6 m_in[194]
port 106 nsew signal input
rlabel metal2 s 166170 219200 166226 220000 6 m_in[195]
port 107 nsew signal input
rlabel metal2 s 166998 219200 167054 220000 6 m_in[196]
port 108 nsew signal input
rlabel metal2 s 167826 219200 167882 220000 6 m_in[197]
port 109 nsew signal input
rlabel metal2 s 168746 219200 168802 220000 6 m_in[198]
port 110 nsew signal input
rlabel metal2 s 169574 219200 169630 220000 6 m_in[199]
port 111 nsew signal input
rlabel metal2 s 17222 219200 17278 220000 6 m_in[19]
port 112 nsew signal input
rlabel metal2 s 2042 219200 2098 220000 6 m_in[1]
port 113 nsew signal input
rlabel metal2 s 170402 219200 170458 220000 6 m_in[200]
port 114 nsew signal input
rlabel metal2 s 171230 219200 171286 220000 6 m_in[201]
port 115 nsew signal input
rlabel metal2 s 172058 219200 172114 220000 6 m_in[202]
port 116 nsew signal input
rlabel metal2 s 172978 219200 173034 220000 6 m_in[203]
port 117 nsew signal input
rlabel metal2 s 173806 219200 173862 220000 6 m_in[204]
port 118 nsew signal input
rlabel metal2 s 174634 219200 174690 220000 6 m_in[205]
port 119 nsew signal input
rlabel metal2 s 175462 219200 175518 220000 6 m_in[206]
port 120 nsew signal input
rlabel metal2 s 176290 219200 176346 220000 6 m_in[207]
port 121 nsew signal input
rlabel metal2 s 177118 219200 177174 220000 6 m_in[208]
port 122 nsew signal input
rlabel metal2 s 178038 219200 178094 220000 6 m_in[209]
port 123 nsew signal input
rlabel metal2 s 18142 219200 18198 220000 6 m_in[20]
port 124 nsew signal input
rlabel metal2 s 178866 219200 178922 220000 6 m_in[210]
port 125 nsew signal input
rlabel metal2 s 179694 219200 179750 220000 6 m_in[211]
port 126 nsew signal input
rlabel metal2 s 180522 219200 180578 220000 6 m_in[212]
port 127 nsew signal input
rlabel metal2 s 181350 219200 181406 220000 6 m_in[213]
port 128 nsew signal input
rlabel metal2 s 182270 219200 182326 220000 6 m_in[214]
port 129 nsew signal input
rlabel metal2 s 183098 219200 183154 220000 6 m_in[215]
port 130 nsew signal input
rlabel metal2 s 183926 219200 183982 220000 6 m_in[216]
port 131 nsew signal input
rlabel metal2 s 184754 219200 184810 220000 6 m_in[217]
port 132 nsew signal input
rlabel metal2 s 185582 219200 185638 220000 6 m_in[218]
port 133 nsew signal input
rlabel metal2 s 186502 219200 186558 220000 6 m_in[219]
port 134 nsew signal input
rlabel metal2 s 18970 219200 19026 220000 6 m_in[21]
port 135 nsew signal input
rlabel metal2 s 187330 219200 187386 220000 6 m_in[220]
port 136 nsew signal input
rlabel metal2 s 188158 219200 188214 220000 6 m_in[221]
port 137 nsew signal input
rlabel metal2 s 188986 219200 189042 220000 6 m_in[222]
port 138 nsew signal input
rlabel metal2 s 189814 219200 189870 220000 6 m_in[223]
port 139 nsew signal input
rlabel metal2 s 190734 219200 190790 220000 6 m_in[224]
port 140 nsew signal input
rlabel metal2 s 191562 219200 191618 220000 6 m_in[225]
port 141 nsew signal input
rlabel metal2 s 192390 219200 192446 220000 6 m_in[226]
port 142 nsew signal input
rlabel metal2 s 193218 219200 193274 220000 6 m_in[227]
port 143 nsew signal input
rlabel metal2 s 194046 219200 194102 220000 6 m_in[228]
port 144 nsew signal input
rlabel metal2 s 194966 219200 195022 220000 6 m_in[229]
port 145 nsew signal input
rlabel metal2 s 19798 219200 19854 220000 6 m_in[22]
port 146 nsew signal input
rlabel metal2 s 195794 219200 195850 220000 6 m_in[230]
port 147 nsew signal input
rlabel metal2 s 196622 219200 196678 220000 6 m_in[231]
port 148 nsew signal input
rlabel metal2 s 197450 219200 197506 220000 6 m_in[232]
port 149 nsew signal input
rlabel metal2 s 198278 219200 198334 220000 6 m_in[233]
port 150 nsew signal input
rlabel metal2 s 199198 219200 199254 220000 6 m_in[234]
port 151 nsew signal input
rlabel metal2 s 200026 219200 200082 220000 6 m_in[235]
port 152 nsew signal input
rlabel metal2 s 200854 219200 200910 220000 6 m_in[236]
port 153 nsew signal input
rlabel metal2 s 201682 219200 201738 220000 6 m_in[237]
port 154 nsew signal input
rlabel metal2 s 202510 219200 202566 220000 6 m_in[238]
port 155 nsew signal input
rlabel metal2 s 203430 219200 203486 220000 6 m_in[239]
port 156 nsew signal input
rlabel metal2 s 20626 219200 20682 220000 6 m_in[23]
port 157 nsew signal input
rlabel metal2 s 204258 219200 204314 220000 6 m_in[240]
port 158 nsew signal input
rlabel metal2 s 205086 219200 205142 220000 6 m_in[241]
port 159 nsew signal input
rlabel metal2 s 205914 219200 205970 220000 6 m_in[242]
port 160 nsew signal input
rlabel metal2 s 206742 219200 206798 220000 6 m_in[243]
port 161 nsew signal input
rlabel metal2 s 207662 219200 207718 220000 6 m_in[244]
port 162 nsew signal input
rlabel metal2 s 208490 219200 208546 220000 6 m_in[245]
port 163 nsew signal input
rlabel metal2 s 209318 219200 209374 220000 6 m_in[246]
port 164 nsew signal input
rlabel metal2 s 210146 219200 210202 220000 6 m_in[247]
port 165 nsew signal input
rlabel metal2 s 210974 219200 211030 220000 6 m_in[248]
port 166 nsew signal input
rlabel metal2 s 211894 219200 211950 220000 6 m_in[249]
port 167 nsew signal input
rlabel metal2 s 21454 219200 21510 220000 6 m_in[24]
port 168 nsew signal input
rlabel metal2 s 212722 219200 212778 220000 6 m_in[250]
port 169 nsew signal input
rlabel metal2 s 213550 219200 213606 220000 6 m_in[251]
port 170 nsew signal input
rlabel metal2 s 214378 219200 214434 220000 6 m_in[252]
port 171 nsew signal input
rlabel metal2 s 215206 219200 215262 220000 6 m_in[253]
port 172 nsew signal input
rlabel metal2 s 216126 219200 216182 220000 6 m_in[254]
port 173 nsew signal input
rlabel metal2 s 216954 219200 217010 220000 6 m_in[255]
port 174 nsew signal input
rlabel metal2 s 217782 219200 217838 220000 6 m_in[256]
port 175 nsew signal input
rlabel metal2 s 218610 219200 218666 220000 6 m_in[257]
port 176 nsew signal input
rlabel metal2 s 219438 219200 219494 220000 6 m_in[258]
port 177 nsew signal input
rlabel metal2 s 22374 219200 22430 220000 6 m_in[25]
port 178 nsew signal input
rlabel metal2 s 23202 219200 23258 220000 6 m_in[26]
port 179 nsew signal input
rlabel metal2 s 24030 219200 24086 220000 6 m_in[27]
port 180 nsew signal input
rlabel metal2 s 24858 219200 24914 220000 6 m_in[28]
port 181 nsew signal input
rlabel metal2 s 25686 219200 25742 220000 6 m_in[29]
port 182 nsew signal input
rlabel metal2 s 2870 219200 2926 220000 6 m_in[2]
port 183 nsew signal input
rlabel metal2 s 26606 219200 26662 220000 6 m_in[30]
port 184 nsew signal input
rlabel metal2 s 27434 219200 27490 220000 6 m_in[31]
port 185 nsew signal input
rlabel metal2 s 28262 219200 28318 220000 6 m_in[32]
port 186 nsew signal input
rlabel metal2 s 29090 219200 29146 220000 6 m_in[33]
port 187 nsew signal input
rlabel metal2 s 29918 219200 29974 220000 6 m_in[34]
port 188 nsew signal input
rlabel metal2 s 30838 219200 30894 220000 6 m_in[35]
port 189 nsew signal input
rlabel metal2 s 31666 219200 31722 220000 6 m_in[36]
port 190 nsew signal input
rlabel metal2 s 32494 219200 32550 220000 6 m_in[37]
port 191 nsew signal input
rlabel metal2 s 33322 219200 33378 220000 6 m_in[38]
port 192 nsew signal input
rlabel metal2 s 34150 219200 34206 220000 6 m_in[39]
port 193 nsew signal input
rlabel metal2 s 3698 219200 3754 220000 6 m_in[3]
port 194 nsew signal input
rlabel metal2 s 35070 219200 35126 220000 6 m_in[40]
port 195 nsew signal input
rlabel metal2 s 35898 219200 35954 220000 6 m_in[41]
port 196 nsew signal input
rlabel metal2 s 36726 219200 36782 220000 6 m_in[42]
port 197 nsew signal input
rlabel metal2 s 37554 219200 37610 220000 6 m_in[43]
port 198 nsew signal input
rlabel metal2 s 38382 219200 38438 220000 6 m_in[44]
port 199 nsew signal input
rlabel metal2 s 39302 219200 39358 220000 6 m_in[45]
port 200 nsew signal input
rlabel metal2 s 40130 219200 40186 220000 6 m_in[46]
port 201 nsew signal input
rlabel metal2 s 40958 219200 41014 220000 6 m_in[47]
port 202 nsew signal input
rlabel metal2 s 41786 219200 41842 220000 6 m_in[48]
port 203 nsew signal input
rlabel metal2 s 42614 219200 42670 220000 6 m_in[49]
port 204 nsew signal input
rlabel metal2 s 4526 219200 4582 220000 6 m_in[4]
port 205 nsew signal input
rlabel metal2 s 43534 219200 43590 220000 6 m_in[50]
port 206 nsew signal input
rlabel metal2 s 44362 219200 44418 220000 6 m_in[51]
port 207 nsew signal input
rlabel metal2 s 45190 219200 45246 220000 6 m_in[52]
port 208 nsew signal input
rlabel metal2 s 46018 219200 46074 220000 6 m_in[53]
port 209 nsew signal input
rlabel metal2 s 46846 219200 46902 220000 6 m_in[54]
port 210 nsew signal input
rlabel metal2 s 47674 219200 47730 220000 6 m_in[55]
port 211 nsew signal input
rlabel metal2 s 48594 219200 48650 220000 6 m_in[56]
port 212 nsew signal input
rlabel metal2 s 49422 219200 49478 220000 6 m_in[57]
port 213 nsew signal input
rlabel metal2 s 50250 219200 50306 220000 6 m_in[58]
port 214 nsew signal input
rlabel metal2 s 51078 219200 51134 220000 6 m_in[59]
port 215 nsew signal input
rlabel metal2 s 5446 219200 5502 220000 6 m_in[5]
port 216 nsew signal input
rlabel metal2 s 51906 219200 51962 220000 6 m_in[60]
port 217 nsew signal input
rlabel metal2 s 52826 219200 52882 220000 6 m_in[61]
port 218 nsew signal input
rlabel metal2 s 53654 219200 53710 220000 6 m_in[62]
port 219 nsew signal input
rlabel metal2 s 54482 219200 54538 220000 6 m_in[63]
port 220 nsew signal input
rlabel metal2 s 55310 219200 55366 220000 6 m_in[64]
port 221 nsew signal input
rlabel metal2 s 56138 219200 56194 220000 6 m_in[65]
port 222 nsew signal input
rlabel metal2 s 57058 219200 57114 220000 6 m_in[66]
port 223 nsew signal input
rlabel metal2 s 57886 219200 57942 220000 6 m_in[67]
port 224 nsew signal input
rlabel metal2 s 58714 219200 58770 220000 6 m_in[68]
port 225 nsew signal input
rlabel metal2 s 59542 219200 59598 220000 6 m_in[69]
port 226 nsew signal input
rlabel metal2 s 6274 219200 6330 220000 6 m_in[6]
port 227 nsew signal input
rlabel metal2 s 60370 219200 60426 220000 6 m_in[70]
port 228 nsew signal input
rlabel metal2 s 61290 219200 61346 220000 6 m_in[71]
port 229 nsew signal input
rlabel metal2 s 62118 219200 62174 220000 6 m_in[72]
port 230 nsew signal input
rlabel metal2 s 62946 219200 63002 220000 6 m_in[73]
port 231 nsew signal input
rlabel metal2 s 63774 219200 63830 220000 6 m_in[74]
port 232 nsew signal input
rlabel metal2 s 64602 219200 64658 220000 6 m_in[75]
port 233 nsew signal input
rlabel metal2 s 65522 219200 65578 220000 6 m_in[76]
port 234 nsew signal input
rlabel metal2 s 66350 219200 66406 220000 6 m_in[77]
port 235 nsew signal input
rlabel metal2 s 67178 219200 67234 220000 6 m_in[78]
port 236 nsew signal input
rlabel metal2 s 68006 219200 68062 220000 6 m_in[79]
port 237 nsew signal input
rlabel metal2 s 7102 219200 7158 220000 6 m_in[7]
port 238 nsew signal input
rlabel metal2 s 68834 219200 68890 220000 6 m_in[80]
port 239 nsew signal input
rlabel metal2 s 69754 219200 69810 220000 6 m_in[81]
port 240 nsew signal input
rlabel metal2 s 70582 219200 70638 220000 6 m_in[82]
port 241 nsew signal input
rlabel metal2 s 71410 219200 71466 220000 6 m_in[83]
port 242 nsew signal input
rlabel metal2 s 72238 219200 72294 220000 6 m_in[84]
port 243 nsew signal input
rlabel metal2 s 73066 219200 73122 220000 6 m_in[85]
port 244 nsew signal input
rlabel metal2 s 73986 219200 74042 220000 6 m_in[86]
port 245 nsew signal input
rlabel metal2 s 74814 219200 74870 220000 6 m_in[87]
port 246 nsew signal input
rlabel metal2 s 75642 219200 75698 220000 6 m_in[88]
port 247 nsew signal input
rlabel metal2 s 76470 219200 76526 220000 6 m_in[89]
port 248 nsew signal input
rlabel metal2 s 7930 219200 7986 220000 6 m_in[8]
port 249 nsew signal input
rlabel metal2 s 77298 219200 77354 220000 6 m_in[90]
port 250 nsew signal input
rlabel metal2 s 78218 219200 78274 220000 6 m_in[91]
port 251 nsew signal input
rlabel metal2 s 79046 219200 79102 220000 6 m_in[92]
port 252 nsew signal input
rlabel metal2 s 79874 219200 79930 220000 6 m_in[93]
port 253 nsew signal input
rlabel metal2 s 80702 219200 80758 220000 6 m_in[94]
port 254 nsew signal input
rlabel metal2 s 81530 219200 81586 220000 6 m_in[95]
port 255 nsew signal input
rlabel metal2 s 82450 219200 82506 220000 6 m_in[96]
port 256 nsew signal input
rlabel metal2 s 83278 219200 83334 220000 6 m_in[97]
port 257 nsew signal input
rlabel metal2 s 84106 219200 84162 220000 6 m_in[98]
port 258 nsew signal input
rlabel metal2 s 84934 219200 84990 220000 6 m_in[99]
port 259 nsew signal input
rlabel metal2 s 8758 219200 8814 220000 6 m_in[9]
port 260 nsew signal input
rlabel metal3 s 219200 824 220000 944 6 m_out[0]
port 261 nsew signal output
rlabel metal3 s 219200 170008 220000 170128 6 m_out[100]
port 262 nsew signal output
rlabel metal3 s 219200 171776 220000 171896 6 m_out[101]
port 263 nsew signal output
rlabel metal3 s 219200 173408 220000 173528 6 m_out[102]
port 264 nsew signal output
rlabel metal3 s 219200 175040 220000 175160 6 m_out[103]
port 265 nsew signal output
rlabel metal3 s 219200 176808 220000 176928 6 m_out[104]
port 266 nsew signal output
rlabel metal3 s 219200 178440 220000 178560 6 m_out[105]
port 267 nsew signal output
rlabel metal3 s 219200 180208 220000 180328 6 m_out[106]
port 268 nsew signal output
rlabel metal3 s 219200 181840 220000 181960 6 m_out[107]
port 269 nsew signal output
rlabel metal3 s 219200 183608 220000 183728 6 m_out[108]
port 270 nsew signal output
rlabel metal3 s 219200 185240 220000 185360 6 m_out[109]
port 271 nsew signal output
rlabel metal3 s 219200 17688 220000 17808 6 m_out[10]
port 272 nsew signal output
rlabel metal3 s 219200 187008 220000 187128 6 m_out[110]
port 273 nsew signal output
rlabel metal3 s 219200 188640 220000 188760 6 m_out[111]
port 274 nsew signal output
rlabel metal3 s 219200 190272 220000 190392 6 m_out[112]
port 275 nsew signal output
rlabel metal3 s 219200 192040 220000 192160 6 m_out[113]
port 276 nsew signal output
rlabel metal3 s 219200 193672 220000 193792 6 m_out[114]
port 277 nsew signal output
rlabel metal3 s 219200 195440 220000 195560 6 m_out[115]
port 278 nsew signal output
rlabel metal3 s 219200 197072 220000 197192 6 m_out[116]
port 279 nsew signal output
rlabel metal3 s 219200 198840 220000 198960 6 m_out[117]
port 280 nsew signal output
rlabel metal3 s 219200 200472 220000 200592 6 m_out[118]
port 281 nsew signal output
rlabel metal3 s 219200 202240 220000 202360 6 m_out[119]
port 282 nsew signal output
rlabel metal3 s 219200 19320 220000 19440 6 m_out[11]
port 283 nsew signal output
rlabel metal3 s 219200 203872 220000 203992 6 m_out[120]
port 284 nsew signal output
rlabel metal3 s 219200 205504 220000 205624 6 m_out[121]
port 285 nsew signal output
rlabel metal3 s 219200 207272 220000 207392 6 m_out[122]
port 286 nsew signal output
rlabel metal3 s 219200 208904 220000 209024 6 m_out[123]
port 287 nsew signal output
rlabel metal3 s 219200 210672 220000 210792 6 m_out[124]
port 288 nsew signal output
rlabel metal3 s 219200 212304 220000 212424 6 m_out[125]
port 289 nsew signal output
rlabel metal3 s 219200 214072 220000 214192 6 m_out[126]
port 290 nsew signal output
rlabel metal3 s 219200 215704 220000 215824 6 m_out[127]
port 291 nsew signal output
rlabel metal3 s 219200 217472 220000 217592 6 m_out[128]
port 292 nsew signal output
rlabel metal3 s 219200 219104 220000 219224 6 m_out[129]
port 293 nsew signal output
rlabel metal3 s 219200 21088 220000 21208 6 m_out[12]
port 294 nsew signal output
rlabel metal3 s 219200 22720 220000 22840 6 m_out[13]
port 295 nsew signal output
rlabel metal3 s 219200 24488 220000 24608 6 m_out[14]
port 296 nsew signal output
rlabel metal3 s 219200 26120 220000 26240 6 m_out[15]
port 297 nsew signal output
rlabel metal3 s 219200 27888 220000 28008 6 m_out[16]
port 298 nsew signal output
rlabel metal3 s 219200 29520 220000 29640 6 m_out[17]
port 299 nsew signal output
rlabel metal3 s 219200 31288 220000 31408 6 m_out[18]
port 300 nsew signal output
rlabel metal3 s 219200 32920 220000 33040 6 m_out[19]
port 301 nsew signal output
rlabel metal3 s 219200 2456 220000 2576 6 m_out[1]
port 302 nsew signal output
rlabel metal3 s 219200 34552 220000 34672 6 m_out[20]
port 303 nsew signal output
rlabel metal3 s 219200 36320 220000 36440 6 m_out[21]
port 304 nsew signal output
rlabel metal3 s 219200 37952 220000 38072 6 m_out[22]
port 305 nsew signal output
rlabel metal3 s 219200 39720 220000 39840 6 m_out[23]
port 306 nsew signal output
rlabel metal3 s 219200 41352 220000 41472 6 m_out[24]
port 307 nsew signal output
rlabel metal3 s 219200 43120 220000 43240 6 m_out[25]
port 308 nsew signal output
rlabel metal3 s 219200 44752 220000 44872 6 m_out[26]
port 309 nsew signal output
rlabel metal3 s 219200 46520 220000 46640 6 m_out[27]
port 310 nsew signal output
rlabel metal3 s 219200 48152 220000 48272 6 m_out[28]
port 311 nsew signal output
rlabel metal3 s 219200 49784 220000 49904 6 m_out[29]
port 312 nsew signal output
rlabel metal3 s 219200 4088 220000 4208 6 m_out[2]
port 313 nsew signal output
rlabel metal3 s 219200 51552 220000 51672 6 m_out[30]
port 314 nsew signal output
rlabel metal3 s 219200 53184 220000 53304 6 m_out[31]
port 315 nsew signal output
rlabel metal3 s 219200 54952 220000 55072 6 m_out[32]
port 316 nsew signal output
rlabel metal3 s 219200 56584 220000 56704 6 m_out[33]
port 317 nsew signal output
rlabel metal3 s 219200 58352 220000 58472 6 m_out[34]
port 318 nsew signal output
rlabel metal3 s 219200 59984 220000 60104 6 m_out[35]
port 319 nsew signal output
rlabel metal3 s 219200 61752 220000 61872 6 m_out[36]
port 320 nsew signal output
rlabel metal3 s 219200 63384 220000 63504 6 m_out[37]
port 321 nsew signal output
rlabel metal3 s 219200 65016 220000 65136 6 m_out[38]
port 322 nsew signal output
rlabel metal3 s 219200 66784 220000 66904 6 m_out[39]
port 323 nsew signal output
rlabel metal3 s 219200 5856 220000 5976 6 m_out[3]
port 324 nsew signal output
rlabel metal3 s 219200 68416 220000 68536 6 m_out[40]
port 325 nsew signal output
rlabel metal3 s 219200 70184 220000 70304 6 m_out[41]
port 326 nsew signal output
rlabel metal3 s 219200 71816 220000 71936 6 m_out[42]
port 327 nsew signal output
rlabel metal3 s 219200 73584 220000 73704 6 m_out[43]
port 328 nsew signal output
rlabel metal3 s 219200 75216 220000 75336 6 m_out[44]
port 329 nsew signal output
rlabel metal3 s 219200 76984 220000 77104 6 m_out[45]
port 330 nsew signal output
rlabel metal3 s 219200 78616 220000 78736 6 m_out[46]
port 331 nsew signal output
rlabel metal3 s 219200 80248 220000 80368 6 m_out[47]
port 332 nsew signal output
rlabel metal3 s 219200 82016 220000 82136 6 m_out[48]
port 333 nsew signal output
rlabel metal3 s 219200 83648 220000 83768 6 m_out[49]
port 334 nsew signal output
rlabel metal3 s 219200 7488 220000 7608 6 m_out[4]
port 335 nsew signal output
rlabel metal3 s 219200 85416 220000 85536 6 m_out[50]
port 336 nsew signal output
rlabel metal3 s 219200 87048 220000 87168 6 m_out[51]
port 337 nsew signal output
rlabel metal3 s 219200 88816 220000 88936 6 m_out[52]
port 338 nsew signal output
rlabel metal3 s 219200 90448 220000 90568 6 m_out[53]
port 339 nsew signal output
rlabel metal3 s 219200 92216 220000 92336 6 m_out[54]
port 340 nsew signal output
rlabel metal3 s 219200 93848 220000 93968 6 m_out[55]
port 341 nsew signal output
rlabel metal3 s 219200 95480 220000 95600 6 m_out[56]
port 342 nsew signal output
rlabel metal3 s 219200 97248 220000 97368 6 m_out[57]
port 343 nsew signal output
rlabel metal3 s 219200 98880 220000 99000 6 m_out[58]
port 344 nsew signal output
rlabel metal3 s 219200 100648 220000 100768 6 m_out[59]
port 345 nsew signal output
rlabel metal3 s 219200 9256 220000 9376 6 m_out[5]
port 346 nsew signal output
rlabel metal3 s 219200 102280 220000 102400 6 m_out[60]
port 347 nsew signal output
rlabel metal3 s 219200 104048 220000 104168 6 m_out[61]
port 348 nsew signal output
rlabel metal3 s 219200 105680 220000 105800 6 m_out[62]
port 349 nsew signal output
rlabel metal3 s 219200 107448 220000 107568 6 m_out[63]
port 350 nsew signal output
rlabel metal3 s 219200 109080 220000 109200 6 m_out[64]
port 351 nsew signal output
rlabel metal3 s 219200 110848 220000 110968 6 m_out[65]
port 352 nsew signal output
rlabel metal3 s 219200 112480 220000 112600 6 m_out[66]
port 353 nsew signal output
rlabel metal3 s 219200 114112 220000 114232 6 m_out[67]
port 354 nsew signal output
rlabel metal3 s 219200 115880 220000 116000 6 m_out[68]
port 355 nsew signal output
rlabel metal3 s 219200 117512 220000 117632 6 m_out[69]
port 356 nsew signal output
rlabel metal3 s 219200 10888 220000 11008 6 m_out[6]
port 357 nsew signal output
rlabel metal3 s 219200 119280 220000 119400 6 m_out[70]
port 358 nsew signal output
rlabel metal3 s 219200 120912 220000 121032 6 m_out[71]
port 359 nsew signal output
rlabel metal3 s 219200 122680 220000 122800 6 m_out[72]
port 360 nsew signal output
rlabel metal3 s 219200 124312 220000 124432 6 m_out[73]
port 361 nsew signal output
rlabel metal3 s 219200 126080 220000 126200 6 m_out[74]
port 362 nsew signal output
rlabel metal3 s 219200 127712 220000 127832 6 m_out[75]
port 363 nsew signal output
rlabel metal3 s 219200 129344 220000 129464 6 m_out[76]
port 364 nsew signal output
rlabel metal3 s 219200 131112 220000 131232 6 m_out[77]
port 365 nsew signal output
rlabel metal3 s 219200 132744 220000 132864 6 m_out[78]
port 366 nsew signal output
rlabel metal3 s 219200 134512 220000 134632 6 m_out[79]
port 367 nsew signal output
rlabel metal3 s 219200 12656 220000 12776 6 m_out[7]
port 368 nsew signal output
rlabel metal3 s 219200 136144 220000 136264 6 m_out[80]
port 369 nsew signal output
rlabel metal3 s 219200 137912 220000 138032 6 m_out[81]
port 370 nsew signal output
rlabel metal3 s 219200 139544 220000 139664 6 m_out[82]
port 371 nsew signal output
rlabel metal3 s 219200 141312 220000 141432 6 m_out[83]
port 372 nsew signal output
rlabel metal3 s 219200 142944 220000 143064 6 m_out[84]
port 373 nsew signal output
rlabel metal3 s 219200 144576 220000 144696 6 m_out[85]
port 374 nsew signal output
rlabel metal3 s 219200 146344 220000 146464 6 m_out[86]
port 375 nsew signal output
rlabel metal3 s 219200 147976 220000 148096 6 m_out[87]
port 376 nsew signal output
rlabel metal3 s 219200 149744 220000 149864 6 m_out[88]
port 377 nsew signal output
rlabel metal3 s 219200 151376 220000 151496 6 m_out[89]
port 378 nsew signal output
rlabel metal3 s 219200 14288 220000 14408 6 m_out[8]
port 379 nsew signal output
rlabel metal3 s 219200 153144 220000 153264 6 m_out[90]
port 380 nsew signal output
rlabel metal3 s 219200 154776 220000 154896 6 m_out[91]
port 381 nsew signal output
rlabel metal3 s 219200 156544 220000 156664 6 m_out[92]
port 382 nsew signal output
rlabel metal3 s 219200 158176 220000 158296 6 m_out[93]
port 383 nsew signal output
rlabel metal3 s 219200 159808 220000 159928 6 m_out[94]
port 384 nsew signal output
rlabel metal3 s 219200 161576 220000 161696 6 m_out[95]
port 385 nsew signal output
rlabel metal3 s 219200 163208 220000 163328 6 m_out[96]
port 386 nsew signal output
rlabel metal3 s 219200 164976 220000 165096 6 m_out[97]
port 387 nsew signal output
rlabel metal3 s 219200 166608 220000 166728 6 m_out[98]
port 388 nsew signal output
rlabel metal3 s 219200 168376 220000 168496 6 m_out[99]
port 389 nsew signal output
rlabel metal3 s 219200 16056 220000 16176 6 m_out[9]
port 390 nsew signal output
rlabel metal4 s 188528 2128 188848 217648 6 vccd1
port 391 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 217648 6 vccd1
port 392 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 217648 6 vccd1
port 393 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 217648 6 vccd1
port 394 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 217648 6 vccd1
port 395 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 217648 6 vccd1
port 396 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 217648 6 vccd1
port 397 nsew power bidirectional
rlabel metal4 s 203888 2128 204208 217648 6 vssd1
port 398 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 217648 6 vssd1
port 399 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 217648 6 vssd1
port 400 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 217648 6 vssd1
port 401 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 217648 6 vssd1
port 402 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 217648 6 vssd1
port 403 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 217648 6 vssd1
port 404 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 220000 220000
string LEFview TRUE
string GDS_FILE /project/openlane/multiply_4/runs/multiply_4/results/magic/multiply_4.gds
string GDS_END 140184930
string GDS_START 411536
<< end >>

